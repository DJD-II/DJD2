    ����          @  ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j����wEj�kB�A~r �x�2��H�"�BДN��á7ڴ �rA7Nm@��):Y�]��/�|��gW�:��Փ]���]�Wd���'��=�a0�a5k��7(��8�t9_����j�sRu�BMM�Dp��{?;b�)�����r/��F������Ό,�]��}��7�I�Ik�H\��Pnd���Y4l?���Y�E���Y�^�c(�w���T�w��>q1��/;� �#'o�Ĭ*�T:�(�^�e��\%Fɯ����[��� ?��`��<�������I̫-��(d:@��C'&é�1D�#)zL�Ԃ�/&F�}
��>o�x�ېy뻑Fi������������_�\����*������~��?~�Hޱ"�yXZC������c��28ג��[�u2W�h�C�bN���*��m��e�%j�k}�"��ȆAK���Si��G#[���>ur�UԠgCF~L���;�i�yqj��^�j�%;�o�hg�#���pn��rË�'#M�^ݘq��fU��|���Q�h�����.~o7��m%��⸞.Z��_�r�����ά���s�sC�������/�6�۩�݅����6�Gl��y5�^a?��-s�(e��f`|����p���3��E�\J�};�ax�����aw��9S?�6��>���2�e�`�C�a�VL���S���5
�GpԂ�eH8*��9�Bʤ�WN��9A�q�u�ɇ:?F&�6G@	�M Ѿ�:�-����]z��̆��%���p��Ѝ�K��{�=���ۻ�2�ҹ�2��h]3$�6��6`�5�Y?U�
�K�ճ�%5���#uk�)��ՄU}��X%���D�y�S��c������H��{D��jl��l��¼�3�7e��
������GUm,��͞O���<�hS��o]��s@�~�ݒ���AR�r��B�'3h"�+ϠFƴ.�bkm�.J�P���\��!�Pw�l��gtM�L��I+�~ɚ5y!~xͥS<[$�l��TW:��'�	S�ÖN��k)�+=���'l�vZ��
h�3��ȿ~�9:�z?[h�ה�xl8�V�QCK⋑�"�z��M�9 �M1jm�}_����2���!�_:����{EF��Af��J3)�{�W�+�c�м����f��O��vJ�$��P�א�]�m�ZR]5 ���8.����*������o��&��ݨ���x�dB��u�}D��?tugcq�)��F�H?OF�
����(L�#�]Fb�� �2��J�ަ�A�i���u
u�uVX�0n̿�W��-��8�́�ݪ�+���)��Cx��vd5TD"B�@�b�ā�{�&G�Js�1HG���TGp5�x.岶o�>��o��*t�`j41�c���hw&ʝ�C�P������;
�+��=�5�.�� 
��d�@���A�)���1��U��w�!T�ς�x>�����/�� �x�N6J3�ÓY����`eo�i7�P�A%��& ��r~ړ��A�@zJA�z�k�rB���9ɧC:zḰ�l:ЕD���aJ2=gE����W���'M�BȠ��H2��!T��P�bڐT��}�8����#Avj?*y�2��=@�T~q8��\��h�윱@���T�M���;ů�m{�v���b)�b�Cf��O.?�Wݲk[y,�2��Iq��\��vM�(� g�1�Y��[�'*���5
��VS��Ȑ�Y��83�jY�a����H�{�ك1=�ڟf�˳�ݻ���G$�B�m�J�N9Q���&w	s=W�$�T�`�m������q��[۠_T�R���č���]X�p�o^�5��3�8��0�[j�wg8Z����������Ş�P���i����}
����\����.''9�]��rĀ1�N��n$���L���;�F��4��B�� 2 �vV5&�* ��N����6K2���^����Yw��&z��JPy��/ƭ�Iy7��OtG�Y�H��~k��b�p3�:)�싗�h��� ھ]���n���+^�>�ȃO�M?s�Q��*�h&�q_�Xq)���r����c�a�wK��΍`)H��Y#�7�We�zWR&١�a��-x��q���S����v�g~�;}�� ;� ��	nsoJ���6.�k�{�Q\P���)�]��}O�z��k�ʇ�2WD[��<TKp���מ��֘P�dr���4曻9�p�&�L`t༘�ez.V_����mK��:~N%��pL��X�iq�\���ya������3���LA����(*�@�}��5�Y����� Cre�L)ū��VEcT�o}T�̝�̃C����ڍ�h!������t���J�Om&��.���-����¸;�]����wL2������G�kF`/�ɂ�_2�j�'�~�d�#� 5Sj�MZ�:�z��9�mN-b��O4�Jk�T�d���V��[ˋV,md�C��ڗ�f�1K��h�n�:���^�T�(��o�4�z��qx/(�B-5��2�x�JK�[p�!�����Ǉ�Һ\����y�8}���Ô����y��L����㐪ß��J� cߌf��)>���[���znQj���"�"�߷�/n�w�z��3)��A�u�d���i�#U�̤�̐���R�w����!aUt��a�Ϫ`�s���o�9������}�\*�:�P7 ������Ӊo�^���%*��)��π{����E��|@���R#1���H�./VHh0�ja�w_H>�֠h9Uv`=.�?�!�8����!u,����|��V�����;��d�������K_�l����FP��;���cs����Pk��Ԕ�|�ݳ��{�P�`�%=�����)��+���	9L�B�Zl�����b���7�X/��p]�NVU�,���a�������#RI*z�M&lMs���̅I��P�}+с8���{�^!�,k�A�H���X~g-�ϐ��Q�o�f�6�ؖ]��O�.G�*�Щ�L�� 4�R�	��[e�.�F�S�,Th�8�X�N7�H��>�ҍCW���}E�ʑv��&=I��b���,E	,qYRl&C<����+�f�ɝ{�ˡa��EB܁����xKƮ��@+{��;Q�S����4a�I�<�����I�]u�BNӠ���9GJJn>��f6d��� ����C���e|�e'(�`J\�T��jԞt�1���Ő!J�;u��3�D�E4�=��mx|RlI���ns��5b����l�^��l0�J$Z��J~�Hj�V��%!c��,�o�ƂD�����Ө�0�1m ZA�%I\I��'	�⾷[�؃�_L��5��ttC�'\{�Odm]�!q��TAY�^0�EE�����w�iXY��st�+w|�v>~�Z��Z�1�_$��]T���B@Td�̣���q�ʣ�+��X�	_�;��wZ�v�^u��y�O��@sl��W|��4E��%e�q�a�x.���>aƅ��<��*zƐ��K>`���}$Y���[;|����iej��+j�I6�����L@�*�IM��C*8����!�8��v��֡F@��2���@ݍE2�}��Z(�"u���cY�͜dk���2������?O�ȇ'��&�(h��6���6џ��V���B���#��$R���.b�X�؅HpکV~N��X[[&�.]y�&^ә��R�ȒY�5�锁f��R��������� ����r1��Q���z�_i�ڬa��x�L�gJR�n��z�[Y^r��>0߸+D ��62�;��I74�mZc����� y<I���?ɺ�֒ʔ-��^�.�'6�<��Ŗ����`A��!.�}Sn�g� �3$\߿�sm�	���Nf��b`�m�nn]ס�!��c����*�CI�f�
� V�<7Y{�a�W��nd��xc���*oJ��TJL����uY�XT�j�{�$ɟ ﶰ�>W~j�j�pqI�2.��*�01���D��Ϗ��|ow7nZ�����$@�^ѷ���8��L����U]�Llk %�N>���Bx]����0�D"���?H��
F���ә�/�-���4�]K��kaa�i��;pY����z�+#"^�Y~�M�)$����;�.��V��j=�������}_F7��i��.������	�rK&h��9X�C$Y<���ÇɌ����%}V�w-�P�c�'U���%4�m�R8�m%by�Y�v��������2!�1g�4��
�C����^�,���)���$����T�(B�	)	2��X{.�6�`B�@U���G��꾥p`���-s�v��]jE��7�8��d�����f��6N^D3���E�z�����c�n�(p|T�"'�R����;���>�Ԟ=3v¯�፻�P�6�B{���z1�Ɉ���AG�Ř{x�r��GH����.�[��F�J�1��W���ش��J��]m�u�ݢ����}�RL�C��D���ݿI5�u�f<(��3�u�u�e����[��U�,N��V���<��6�w��^Y�;�z��z)	��`u��X�i(�<�������5�Q �#̼�1.zo�ˌ%�S��$^3ҵa����*%$AcV�㈓h�l�ڶ�����D���RB��Ca�f�mwx������fzӣ Þ�
h)&���Ic�a�A! ᖟ�س41�@�;�ʩ�|j2.�6�� �e�6gir������ѩ�56nJ�![%Z���u�*�8�2LO�W�Z�wIE��4���߲��J:h^���ʑ;��;��7��K�R��:���8��fU��f��]��C�ɪ�5\w.��r(1FJ���`�e0�R舋sAƟ@���l��?�GrO�v�tp���c�g��
�:��4A����چ���M씃A�cA��=}X��R6l�3:�"k�\�T�=�N!���U���� �Rɓe���cEGO��D��l����ӛ����4CE�����,�Z�.m���U�x���+e�8��gS/ޏ9���y˛��aPg �g���u8C����)�S���I�v���:�d�V8Z����&��/��G_"j<���%��Z��K��8�V�T�ع;B6��>6�k�u�T�@��!�`8oJ�ݽq���������T��'>c����U�r/���FWZ-��?H��W���c���/�y_R�B��ӆ��P�\d���av��AF��?"/��W��gg�x�>�	�曱�_�]Y@��\�<?&���B��!{}"�=���ܺ�؉��e6ۡ�pR[����Lw�-�΀M�Eϒ��u��%�YQP09�Å'�\_.y�)�ɥx~��?��D ��s#��3Ւ�WY�,0f5���\�jD_1=2�P��h�
c��.��͖�:ƴ5���@�+ v�f��*e5��zrJ��axw��݂��<��H�.l,N����$dx�c����x*ԟ�����Vv�q�����q�i��n�S!�Ŝ`e��;)�E�׼��+�m:b��ÄydI�W��H�{�B����~��;ã}h%�m�:��G�W�b����E������MD�{<c�[�U��hס�)��b�a~�vؐ���0JH�/�p�!w�|���
R8��EL��Up�␳�u�Q��-�ZJ�������؊��{�׮H΅�����7H��cOä��g_͓*_��
��{D!��L���vrC���>dW:ڎwQ��N.@�,�}�H�o}����</���!��H��W� ��.���������J��O-Y�.�6�����\��y�<����r�ܙ�Ļ�ʎ�<�����޿��	��&�@/�Wl�1��#������"���s*w��� J"���P�Lsl3;�jL����o�.��.������2K�x����Ͳ�����!~G��p�J��%B���ɐ	B'�ׇ������,����bZN��yո�� λ�j��5m��'rU��^�����z�֐? g����(�7��E�!�^4���f�hI��+���pJ�yDk{&3��M����"!S�����мf�B	��C��ә�<U�2�A���lFܸ�cg�Q?�J���9�	���bx쾮�����*̶�x����BI��4��u�w�#���=2��[}X.��(�'W�t�9?�U���f��{�ا� =US!�Z�#�,��=���˕J�/�%�x�\�p���՜=i��.Bc#��R>����<z�z��r�H ��I GG#�}��^A�w.8����ɐ��ӝ�z��3�l�(���z;�z^�8̂�I��!A
oх�uڲ�|-���B�Dl�%�X�cF��|�q����������)gA��]z������d����=�ty�m̈3N��Nyd��A�����\ �qԗ�#��~>-ܬu�O�o;ЭZnQ�zʅ4� ��� $~5ݣw��~h�v-ɟ��q�2��+@�@G�0��ٷT56"���t �`uX`;���y����L�4=�%� r���`�?�{���޻Y��Z.ůu,t���@��LPQ��s)���c� �����9�6w��.���+��ݰI*��]x����֣�w�J��M>;�,TN��C08��?�XQ$~Q��8w���p��}��sAQ��t]5��0��_\�S6"ơe��%� ���޹�4k�N��=�g?k�s�<�a��7�:x:�r�t	g����]�gG�.3�A�Y�ֽ6��+� �}�=�ڎY-��gQ�����0�q�tU*���J�EA���Y��E�+A妚���oR,.%��ж�{��V�L=?��-!t����v��&d�sxj��瞿�S-RI,lʃ�kx��tQ�UHju�g��|�M*��W�|��P��%�v��Qn~*P���<J>M���z�����a�� �]��?���:XX���g��<�+mk6V�"���+�:\+K+�/�Q�c���ޚ-�Ĩ��=oq����u(��:��i�I�*�[c�^���4�Zuw��o0�\V��8�������*�͒/�e��GWI�G���˝�L��w��P��/e#�)S��ԽW��_���e�֚�l�sd��2�b'��藯۰�#�r8��rsH�����]KГ���M�	-Di�4�����[R)V���TCy�:�k[��?q������>@Nf p�ܛ�w#����籿�2Í�~����}.[˃���B��c"w�4b�
(ǁ�r$���
+���(�*o{C��߷��u6K�i���N|����D�r�d�&¢�㠔�1�v�b��A��g�E��C���L��tX�Dy��o�.�q���|.��G6 ���0��y�,f���<��Q�<��XA6��DW�3�0��r@W��g�ʹ�����2׹e�w����i+0<ii�yI;]��/�^�h	O��H�J|4om �
כ^*o"�a�4�'�B�M�E��1aE<�~w=�\�6��_V�,ZL�E�}]��!8
������݆"s�t@Шr񭙒�ZDÿ@��F3�R,����Y���ˍ��+��ѹ�'��:��B6D'i�t�Ů�p�g�E��c-�;���~c�E�=����6�����s]S�X�I;��.�!��O���K5w��q�y��jQj�E���lG T��M���Hi4������y_��#�=�q��Q\��F�A>G� ]���uւA�e����:����d$g��~���U�Z((:8a�P\�{B���i;����΄fZ�z=�A��v���}Y��
    ����          �  ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j����wEj�kB�A~r �x�2��H�"�BДN��á7ڴ �rA7Nm@��):Y�]��/�|��gW�:��Փ]���]�Wd���'��=�a0�a5k��7(��8�t9_����j�sRu�BMM�Dp��{?;b�)�����r/��F������Ό,�]��}��7�I�Ik�H\��Pnd���Y4l?���Y�E���Y�^�c(�w���T�w��>q1��/;� �#'o�Ĭ*�T:�(�^�e��\%Fɯ����[��� ?��`��<�������I̫-��(d:@��C'&é�1D�#)zL�Ԃ�/&F�}
��>o�x��.����}����mW@�=����	h��EE���դ��H��"ّ�<5It·�9�U�s��T���$�#=�3ۤ��/�ʆ�����`�UO,�ğ������K[�i��C7��A
{�Ƥ��?� K������Ƃ�z�� ���"Q�&��QTa���d�.$6r�+��$c(�)$�����g�H����ޏd� ���y:E���}�O+�Q��X��;NhԹ���tƎh*�88�D���H�.���K���<z
lvmG,e�����7=��5鈮g�C�c;�O�,���=���2� �`��J�9���ȝǫ���Z�Hl�����v�ģՂ�O����lbg��E5E�����e"���P&���g��W��݇��,Jٔ�78�8m����� G�Wt��[^��� W�b#u#z��׈3�g�掵+ӻuQ������_�~��sV�'��� �\e$8#��c����f'iG
��l�����u�e6U��Лw�����9X���l���y�!����+���]��/휠t����:F{I|rX�� G#WP�X|^f/���������ir~vRZS2�����>�_&}�<{���JV��V��{~�:ƫ��t�!�qd�fck��<yh�l����XB|(�q����糛 ��[@��M��� [�':0i(ť�X�o�Q����Q��2P3�\����s�i-@5�9
,]�IrP,����W�����>�T�h�v�CK�L�o?U�����A�P���A�O&����s4�l��W�!� ��b-�ث�����B�T@��yB�ze8)ne��zF҉�M!�E!�<"�{��J4�FCm1�k��`U& ×4!^~�ળb�&�-b���*ʢ$N�k:���u��[�K��6C}}�����y˦�ֺ[�F)��$��1Gn�åα��T(^pT��b52�3������S�����@����'X/�<�:x�k2�D�z�k�'��\̥R��(��ZS]���ں��p�Vxc�U=�~U8<0�k�pF����Ո��/�q�lo��=[%2��V^���0��:d�	Ȇ+%�/�j������,2�w�@�!v��ϫ���5����������p�������J�*��N�H�CZ��TUR/�%�`Rp/���I�J�|\���*�4Ϧ�=\(���>{3`ѼpuAZ��3��T��E:2�4l�wwP�����I@�1S����b��V�y�2ᡭ�Ѵe�%��b%I�X({�~"� ��T?`���ֵn�l� ���Cu�ٶ�ڎ2k��Zy���o��8�����z�'{u\���8�u
-|��	���w�<�����{]�!�|ێ8�t��l��@�ĕɵ~y0�",;fjq|N�����Z.�ġ5��{��N.�>E'�)����P���ޕz��R��m�.{J��T����$c}��<��X{v"G��<��Nm�E��{L���8�t����c��ńsJ�A��$�A�U��������s��#o�>��}xG�N���'�o!��R�������t�]b��.8 �����	�y�\�Oc����3)m�0N�Ź��b��!�,���`�L{��QN0�4������ �D�֣q9SpЏ��2o���ݹH�>��ȗ�TL�pJ,�}�����VC��P�Qg�sw���^�9���Q+�QԤ�r��AڝD_�S@H �A����<$	2qA})K��\�rus��Gm�xE�>m_��(2Y�9�gr����A
���ht:��u�ЊX2�ߒ[-S��ף��LC/4vd�01�E�ˣ?̇��8b��Js%�m�+�?޻���T�Y��B�M��)?���3K�|D�Q���P\q7vdM��O�0x `���Uk�nU�N����p�Etd����D	���n�
���A� K�Vp�t�:�KV����OQ�����Ց��-��k����׿$�F���qȋe��r���y��5?�QX�S�+fu+��ήI�*��)�N�;cgU�8 �}~y�M���)GL`�E���u2�@�Z����3�.��F�ͳh�3 ~2��i�m�x��sm��zw^e��Oʪ���A���w��@�E�_u/:����[fs�����Toj�IW�d��n=���E��zgؔ�pӨ�+�h;UJ��^�'��A��Q��*" ��E��t�s<lᆱ4 �wmJp ��=G�R|˾5#ͯ�j�a N5�Ư�K5�L���N'�Kk�iu5}�}:�>)�C��	��۷�����YC9�= �F_ބ�5�l@��� XJ*�sL��*�neW�U-1tƮS�C�I�	��B�iPC����1J=-�n�|^s7Ϧ��9���J�,sz�hMf��xf&W;��y���֙����0��-ѿ;Z}UJ��K����*r���.��/��c��U��:=����5�j�GyZݟ)��'�)lXNWəe�0�3K����=;vu$p]t���};}�>^�!>�
���$��'!m�d����>�&��Q�JI���Yye�ko�ƪj�<������s-�*Q�te�7�xjxl����BAԎd-<�=B>k04���u 4Ȓ�m5��[N��_(�<8w2Y�3��Z�W/�h�D�ѽ.-@��bޭ|��n�̈��S����d�S|�-ʝk��c��T�X��oCϙ��7��A��v4뻱��M�f� ;8Q�q]��#��-�#]4��'��hWHqE�z�g�4���Y�i gxjP���1�������0i�P}L���zQ{��v�]⦣D��S	�T�nʐ�S��c�ə{,}��.<m��޻���f�vz��m��<Y�T�ₛ��_�iCQ��%��]��m@ߜ#4��"�l$�� �Qƃ|8橁!^�Y�T��6��a�&���������[��+��,#�C���\�|��$Ӳ���u��Pк��۬��G���R�d�P��>��Br�]F���ƹ�.��=���O�w�������j˝�ׁWO4�� �s�Y�Y��@��H�d��`L�ˊ����:5�'�er�e2!z�r^�c����+�R�%�_���-��m����!ae=��v��@�b�)�(PV2&����� ������Wv���j�5��	�Kwn޾��zh��%5z�ۅ2(�
��K����+�]yJ���5�2giT�>�\�3���ÿ�`���x���1ԾCF@n2q&3�~ 1{|�����
5��	�u&�	�:F���������x�r�J�dEӤ���g��>c�1���
5Y��.�ԁG�P
�4���z͒�Dpr*��H{ ��jcZ4��+ C&c[s��Q��/�0�cąAXM��*;��$��4V���oMC�#�m�4�<?���^�ͅS������S�.�ܒ}�!bq��
�	9�z�x��0��W�_G�j�|7U΂iQ��}��n�4L%(�'�q�-!M1j�^�x��9Ĭ�$�����`��i��*���GO}}�'#�"�2K�4R�`q��$��t4>���ޗ2=A�d�ֺ���D�{@��y35�n�\��UWN�ӟC�V]�¡��Br7gJ=.����9TrRP���=|y�]-Rc���>C_!*��7~��b	�GU�!;=/�Ͻ��>�-��1��h�$V���@�6!�]����m�������'�a�Qobb�J����&���o���WIK �8>�x��S�\����+|<�V��T�/�~ �#kS�a�IWt�a������[s�e'��yO�pg ﳢ�ˌw�:�T�,L�l# �^R�s0F�������W��T���)G)��8�R�QOj����>kd�n����]K�2��/��qJ4�	������6[�,O����t�/kh��V��;(w��7P�n+��w���]��ុ�����%l3���c\���Zgƕ��Ki��/5=�$Wq����yJ�cʓ�f1�B����,a%�*�Yn͝[�D��H�
(���'�ض��L�Y��7��2�I�(�p}���?�s;*��8���D��,��p�%�>4T��o}M��$m��Nv�;����E��r�J��.��i=~y�틭_���߀��R�u zo�}}� ����d��)�ߒ���U���9j�aD��lQ]�+�S�V0b�p�o#Z�Ɯ,2������ �C�e��;�Q��O;�$�x�%-�F�j8ew��PC751x�v�C�9�B�F�E������)|	':E��d^�[q��ٔly�/q��N�<쫕b�2��ޞ����+RV�6
]���eo]���a
� 2��<�F�4��Z��[ ��O�x����-�J[��
~���Ow� �5z���94G���_��q=+���hfrǧ��k���X�GT��	�3��l�ոĀ�W�~j=�5���
ے��z�y]Z����S��y�E���K�c�S,��4�����d=a��,�|'}�G"���5���Q�,����o�5^��v<�i���CR����iv��lH��W#���:	�8���dزn`���(�m�?sǑ���5�̳���[(Wv������}�2%h��6�?Ja�������3zHu�Zqw�o\���_�#�[��?�d-�lWPP<J�_�zJKx�~
㾪6��Q~  MK��l5��4���R�����bJ��kC#7�Q��l�Ӥ�^!!�-׮+��	���K��J��_�����6P:6���f���k�<?�[���{��L�C�!�,C�W�'Uv�'�ʘ��� 7Z45��h�o��ɶ��/0�6"y��.�8���ʄ�e+緞�¹�h]թ���0!��s���9/C}��htwüUEߕe)�h��:?ʏ�`mƢ����7���\65oZff?.�jx\������lJ}��u�Dj�d�N�:r��w�ѱ�a���u�=t���/d�����%Ǥ;�ф:�����Z��w�Ӱd��L���7����c������W��\��Z�����ܔi^��CȒ�3�+�t���]��]0:�
��W�gC-�_]g
���K�c���^Ta���Άo���n���`��^k!&k��#9߳C�\Z֌c��V��[��S&�<�Q����<�7X�
4��ؿB�P�ڹ��g^Ļ�X�E(��kBc�����!���a��O�#���U�N�Q^�B7��xK�Kj�D�[�սh��X�K`��in5G�9�؊�>��Y{�G_�\�IWL��c���S,�QɀȤ��;7���r���VC�|5p��Q��8-j��y�X�.C nd1�rp@x���Hz�f�c)LA�v����7�gE���@�5����`�F�dY�� 4>C�4 �VYK��A��k�9�+?��Z����#+x���~A.!%"�x���lu�T~o�=X��"5@��9�m��!�:F��u�i���!x��f۵s�jtWmD�� }\�1L��!e��� ��n�.�\�81"�7����ܳ�>>��%Et�夦?�
{��ɱ�.گ�������P�hjAn�Oj_�S��A���}��f���.��
��b�b�z�w2�
]H��ʈ���ԟ����RTa�ɚ���������=pBU΄�G�_BޗWۦ�C&]���*�G6�@��ޜ1�0�#
	��,N��/K�D:?�=�6?���'��s`��y���DҎ�[H;jۦ�i�6�fp[���M�ȉ���c�C�ё�i��%.Յ�W��uu����V�>Q���Mt���0��v��}\" ��;�8��D?i��K��� �
*-?e��8ۗ{ܹMH��]�j�t:lVU�r=ˮ�hX��j�հ陜=�����B����E<�V�b�?_�24��~�:��l�E�]�y!P�pK�+�Hn~��R����v���j�Hj}���\�oQ��q���	�	~�._0�B����W��Pٛ���5~����V�^@�e��jpW�^�]���V3�oa�`=@[���!�ʓ8'�P��sc`Z�����M;	�=�A9��o�ͳ,id˨߼��F�64F�z�"��W)�3�PS��P]�#�qkm��ސm��Fr��|�S�FԳiG|=s�B�w��5\�̡�L�L�I�q��б�P��m &��}��Vla��q�Nj�{9���BV|Ď�8Y�6lN�1U�{�R�-B��7����P6�S�:�����t��	/�<-:R0��P� o�˂�N��S���'�(@U�����1X{�\�fLnCO���f����6�����hM�+�����Փ����ee���J�9I��hb\�ݥԏ�1<��U��K���p���E�,`R˿7`�q��8��u��!�I���Ё V}u��{bxU=`��Chd�Lcrr�K&p�B6�J`{ֲ:��}���Χ?�8
 �-����8���������fH�P��.�J�yl�6���=�Hx	,sW�C�� ��/�	=�� �!y��� �8<:�a	<nޏ��x̭^��%�/��N���o�� ���n�������y��e�-��@i�X����c�*���L )�1����	�h+�������!��<�y�h0ߡ)7�C�9I>�o�`u����_�9�z7>�<�����22�+?n��k��!�ӨD&���.�z;�'�)���^J��cBN�$$�Z7[$���I���f�(��^V ��*�縪3]	f�w�H]���;�cHq������ώ�sH�u�b@��|G���hԳƢ*Ojp@󁵸a���� �Xh
 ��L��}{���R.�,�Dz�v�(�i�c�vP��A�o��a���[�\n=РB��Q��UU2I��g��@9��'��qX|T�1�����(�{jT%����h:x((��$�}k���Сt�o�"`��LL�yt��>kG�7\����PSRK� &;Ϧ0���քΊ/�X�����M��5/J���
�)v�Sm�(b�؀ ��*A���D6�v�����_����^�>�|:
/m X��%��^��CH �x
[+��-	�e!(1R8S ��T[p7e�Ӳ�@2�3��gi<���w��0�c���Wu�Fy��I�)v�h6Xs�[�Я�R���d�{��#�G��Eﱆ�Ҿ�d?X���?�as���G��4����s�S)���yo$����f����+?��E�&�	����?@�k�@�'����6T(�Aى��Cѓ��fC��%�A")t�X5z7��v;�/���6�-�`q�"PMjV;j_9^��*���Ԩ������x�'�d��T�ڣ�T)Y�OY�����[Z\E�/����rn��&�J��9y� ���7aS�}�����.��.�k�`���,���x��(���*4�U���U��������J��fc��bQno��m�wt�
    ����              ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j����wEj�kB�A~r �x�2��H�"�BДN��á7ڴ �rA7Nm@��):Y�]��/�|��gW�:��Փ]���]�Wd���'��=�a0�a5k��7(��8�t9_����j�sRu�BMM�Dp��{?;b�)�����r/��F������Ό,�]��}��7�I�Ik�H\��Pnd���Y4l?���Y�E���Y�^�c(�w���T�w��>q1��/;� �#'o�Ĭ*�T:�(�^�e��\%Fɯ����[��� ?��`��<�������I̫-��(d:@��C'&é�1D�#)zL�Ԃ�/&F�}
��>o�x��&�ٖ��P| @�$ܕ_�ܘ��r(�n�ٖ�����Δ��O�6*�B��^�,}�Y�U�$eg Z�C�Ys=ܯ+��r��2��T0]2o��i��
�(d�e��J���W���C�lR&��.�Kv6����_�bY�|�� *��d��/���U[��+��p���tsg�3S��*s�c�R
}��}Y�G+ ���Z�S���+�bjN�Y�$W,�����	Ԭ�2��V��{�e3�h���~���#Q�3�Wj�|��H��`�1��u�j:~E�m/g8H����S���Q��(m��%t�H�� ?��������av5�>.:_^�ⳡ��0�^DaCZ�T��R&��B�Lj���j3MU�P���W7��P|��]4>��]��5�|1<G��ͧ"I�|�^|<����0\�}m?��dIg�4�wz a�[1���)Wn�'5�]��n!��h_�K{��U��{�1iLp�զЋ2w�R��0TB�Tm� �����3�ӭb��iBb�,�}�5J�V�'�S�l⃧����!��*ُ!��{���ÿ�[�.�n��˓з�H�k�s��R�H�Eߢ��M�sSP@�G �âi~/SZ�,����?P)0�KO�
���3'����{PΣ�˾�������V�?���L�jsͪ��x`[�c��N�6�� E"�n%a��<킔y�������[���z����J�J�8r�/��c�B�K�%�����N�m�A������P�u1񃱗JQ��Gv���U`�e(u."8��ۚG��7�c�@�92����Cu�7Ը�"��p�Wm����]J�,��W���)ܶD��#�
P�U�a}�{���A(�Ɠ���W�"�U-�z͊n�S�K~W�hM���J�0��]��e���{��"�(��i�M�J�0����㥱m�\=Q���lBT��=�&3�nn9��4�Ud�ms����:�����ǘL�U��ƚ}�Z�P�|~������M0�R���C�A���ߦ�=�f�E��c/X��0���>�s���`�@J��KD��{vi	�ʼp�ӒWȏقd��eIr��B,����6�"leXk(E��.IC�k֭�mi��`�i�Y�;g�LA��h�ۜf�v��늻L0�b��[#퉾��	(dyْ8����"�2л��%���y���W*� 8���QF.��)lr ������n�-���7!T8����7c:a>���oh����Ө@��B��s`6l+�غ)^���#ڏ<
����������f,/�f�D?c��K_|Q&�儔|���H����0���ř�BÎ�'��e�B6DA<9 �p7�X���l���+/��"�y�]:�=@�����w}x�m1i�BMZ���(6�l�
,t?�W���=O]Y�;��uدF���R���N�5��+�W3�r�},ZF����> s���~K]=rk�*���K����ʆ�^w|�����2���-���`�uz��9������x��O,I:$t��n�I鵟޻�0��_�u��)��l{����g��kn��<95�A�=#7#��+��m��@j��$G[8QTB�5ގ����
�B���1��I��j�߀�8�8��2�y��A¸��5�X��	����8 &���F��yT�i"�Vڳ���0�d�H�Gl��e�a�d�W��yͺ\Ղ�Ѹ߮�8r�{Z��cӨo���k�L�J8&�P5�&ݔ�o>ߝ�|�~ڌ�A�m��)a��׵Ke%�����5�]/\�ܐ��x񒖥׼«�hPuq̽�-��7�4F6�����Wg�ߚz���w�N9Y\���������*0�_D�z���ޓ��x�?ɒ�@�m�_2���\>�w����	�L3t���P�M��y[��[@%�uc y�s!�<[�۞��pXN�cHi��=c[6Y��P�þ:=� F��`��th6�Or`�}ʊY*��p;@1��Z�.�ş��z=7M�v;e�����3o�����^y���+oN��`/��O�`�Mƴ���L ��ƾ�{�M���A�$pؔ5�����u8G#C���(��m�s:|x��=[���_��"�c���B����mhW4��K�9�Pk��k�/*r�4�)�͞�r�~/ǰ&J���0�hk���Ak
��G�+��z�������zL�L#��%K�K׼����/Y.�D������`�km_k����e��M&,T?X�+l6� �"��{~�ǰ���8���č��qV�.v���Н��l�c��R�����\>ܼzV��Ȯ���Ɓӗ���#��%��^{n�r��n�2d��q��7"b�I�s��y�M�<Z?���ĔQ�b$s!��ͧ�r,7o۩k������9�ɃT�^��Y��`��7�| 1�����3�V���X�"�]�A�]ŘBV�)��*n׵�5�}����W�l1iЉ\���6<G����hui��P�(1]�A��O�c~xe��۾Gr~y�:-e=��9��[m�%b��Q�:i����+�uKl	�&��@��~`y�~��7K�Y�ĮY*�����p}7
�MV�$�������6uC���������5!擰[)�E�#�9(h�C9{�2�5�W�^�{rf+�w�M�5��B�o��!�e�ފ�B�暻�J�h���}ð����G=Cv�U�E"�|�xC8;�^%hXA���G/���W�3�6����0�(��U	�+or�צ�T`'_��:�	U���@#����+B�hk�c�9���	\�͠ɬmP/b�s.t���	�vlr<-��椺�)���L4��A%�Eo(݈�1�QI'Z��κ1�� 1vC�E��f�6 �F�
Ӿ�ax9��w��ꉃ��սr�,M~|Y�h�9�g���z�/��:��m�y�����Af�-B��l���e����������b�-ҧ';U��5���YAn:1N�H��|zE��#1����Sk<�@�w��`�]V��:z-�Cof��`�jטe�{�=������?��?x��ymk�x$t ���c�n���n�n����\}څ�� 4��������Z	�f��K�����m̋�{c�&���b:�|E��-C��Ͷ&f�).�]��]�/��R�e�^_����OԄx��J�ںA���C؟ό�D�ݑSf1R�s*�0�g�l_J��-���a�8C [H���9=|G�:�+Z-�z���O���r"��k�'���M��@G|���sx"H�bБ:6-n�����6}$%~o�!н�Y���X+[���7R%�W@������!��lȕ�NxtD�u
U�W�AF�q�vvb%���> "�i��<�B[�A>i�'���gTK����*�#u�Y>�lV����0�/饗	�9�㚞y��qb�e���*�uT�nw�ƛbc���C`�0��Q�+�|�quE��--O3�Gk5�b����l�F�kU���2n� u8���9J|�R�KW���`����������D�4@��]�vOٜ�eT��+!�U���j�M�<Gܧ�\ܔ躉!�@����q�kR�w�������J�[z�LZِc���R��A���v��A�+��z��u�bh�l�܌��⟾�ң5����<���V׶.��h�\���O�AVV12��2������`0��s�m,M�J�>n%�Se\�7���c�Z�mRj�5�Mv�F�g1L�g�Ȯ��r�U�;=,_"��� ��D�w�晉W�߾���{F�^�,"�v�G"�`WH��xALu��]�	�[�k�%~�No~%y���&�F�(A
����kZz���z~�7~�c����h4��_FUvuPy3ن�r�v�����|i�}��U-��'��\!�N����o��!ڥ����gq�����tJ�!���?Z�AVN�5��{!3����[Ӳl����H��NJ(����sl#2���E�����٠�AVQ����O��A��b�lh����_�{��r���Y�8#5��}�DM�&.����^?��L�T��iF1k�\��WQW'�M��6���P2���O�꼠�`������ �Ъ4��p6&Z���(| Q?z�����5[/kW�v�&��1����^�*��s� �C9-����lm~2W���:.?H�gq&�K�.r��wڀq���BG���	�ځ�I@������3zy�%����:�{:	Z�ͬ�����\U�t��}�k���[��P������!eIPD��]�SЖZ�By�c���OA�@���ZD1�>��.1T�a��LtkR�^'G��^����G�W@?�`t
������.�����(������`p>	���|��@����5�^i��R62����j�H�{��̥�u� ev"��H{{RC�Y	Q5��TVd��a���ۃO�7g�C�����#�tv/=�.�+j�u�m���ڌ�[�[��D�:ȩ�#���tf��) u5G���fߗT��oC�f/�=#�>ΧX�bld?\*7��������n�����Cxo�H�qk�C8`;I�v�g��p��$@=N��^���!}����.ŗ����Z�0�?0^�Zms�S'�*J%�u�U�}9���hHtr�r��U�héi��w�	a���Q��v4I�S��t2LW�ߏ��
r���-ݛ�0o}NKqJ��pZi��H)��j��4��_�F��/����'W.�ۉ��:���Ȩn�t5pu���˂CU�ϕ��d���}�#9�]�2�6�]c� ��P8�����cG�ߕ5, �I\��~f�?� ��3q =���Od|���+�����g�S�F�0��	r��Kʐ�v �}�����@�`��o�ZN��a�p�b�"�]5���}��O\!5óUր�4콧}8��vȃ�;=���|�����H�&} �����QG�)�/"�7<�=�`?K�L?��ɬ���!����;��Dn38���Vh�jǲ(��ܔ���|�v���ߡ�e/b�*�5y�£҃�)��o:��e�\+��<�����9���x杜���`4�K�C!�4vm����P�O9
�R��&��5�)z*1�68xH��#��M���~��a<A�s�# O�WWf�j��Ш�ty�K~k�XV�l
�^����*E�4���)�"^��-��p��v8����x��&��W�O�:yA�3M��/�\�tst���j]�W1&�ND�*�L��d�N8�����i9��CH���O�,�lH<yƚל��?�`�n������X%x���}��:�&j�"�M@n�*��ߒ��순W<B���-�:;�-�:0�s�ۤ�<G
�я�fA��O���� Ǒ;9�TXi�'�}6n�J2cHA�h��4�o*�o�5w�G���t�v�S F�Y��`�{�k��iD��
�n�Y���;��� i].r���4�G���"P	鯀d��5E�c�$�7�`?^��ü�����眤X~	25��)3Qv!˂�8���.�=�v�Yݤ�Xe�	Z~�X��g�V�4@j�pNM�A���UmŎ&ߨ일�:���=U�����L�$��y%�.����vcQ��e�b�y�^�����u	NcU�H }�1J��M�yo��?�=�����d��4��Uf�_�ȑF����/H,3�FR������{�+es�YV�G���D帣%�!�S	ś&���9�CI�!!�e+�$dr������Տ��"S��&�X@�ܳդa�#�;�~B��~:�����E.��*VǡV~9�>�F��k�zO3��\ю��fJ)Fì������O!4̣,�nn};z�Ĵ�{{9n�������`MSݺ��s�R�]�c���_LrT�t��8x�	""rx��[��/K�:���m	x-��R�Jǚ=;��Qk�+2/�ݫ:�[J&����J�i[��+6�q�}��� r���O�)��͹Ҡd�-`�s�F�����+�W�Do�u/P<�*�G�O1����Y8��oj9ç"�xC�>�ϳ��a~bۦ���glR6��&����o�[�d 5���+�q�����K_G�X�s�g���U�q��]���*�E"�,[�][d&����H&c)�DUт�h	W������AO�:��D���X���8�ۼ��<go|�ZJ�~�s�!��]���!a�n���+v�CzH��.v�e�������tJ-���$b�d������f��7�hD�r~'��ݧ�_����Q����;�f�Rҟ����Ԩ%s�?��E�uQ��c5�E�%�oE6�1R��Ŧu�����+\%�އ�O�+s���9�����u�fin|R*)>n��?]�
L8���&zK+�W��ӺJP�0i����tA ������Feg���5!~R�5ۖ�S��G����E���p�U�4��3�d�:ْBZ�wT
tśS�P��+�
ڝ��d��� �lnz�6>7�i]��^��ĭ�79�Ȯ�S���7����nj..-����RW�<a�}�ν)����l5_l7Y�qC�W�F'�TE&�Ӓ���U*v�����'9�Ģ:�O��	����= "@�ql��PZş���nn�x��}�����p�K�n�PX>�!�iL:��H���4:cWh�k������,/��1=��#��~�k�77��Ï��L�V��D����&ۊ)F݁M���i��k�%�I`I#0���(:�U�S3X,{~��!`����u4^ק�)X)f�o��W���:IdU:7����//�{0��Y�r�l�g�|�ca�:w�6=icb�a$K6*Sc���;���
�Ēv(5 ��I�M�3������C+��7]�NX!��qnb>]pZȘ��>e����\����F���D�?��ԣ�<�	1�E2)�,�**=&�g�	-t$=�A�lb��,�2�!�޶�M�.�������}��p�wN���7�֯O��g.�=�M��k�jgC����m�Z�``�@Fg	*��Ex��4�ڡ�3�P��o�ٴ!Y���:�mu[s�4�̼c�����0���:��s|�b8��g͸T��[$jx�l����
%�>UX`��dC�@��[�����H��ɗ��	!^;����R�]Ry�ȨK)6���,4������}Y�>_�YB���!�w���HX\X>4I��+G��6��R��~f+n��s���"�	������L�(�j��k7�/�!�2��)���O�g�j��7�~���o���1����3G��A&��U��/E�k]$9�\���K��J���f��	�-ד�
O[�Q[I]�Vw��k,�ߩx�i����ov׃��6,1DMKI�� 7����CGo��2���K~�Gy-�,�����H�X����Q��k���ݢPd�������c�D� ��B�&'i�0m}�PgS��Ջ��\��N� �BO�y���[1��:�"3 ���8��s�Đ�EW�>�r`$�J-�T�1>fhs�F�t3D%��˓����XB�B�"���x8�W�4*��=�.���8�;�+�A6�� 
>�8�� H�\�x�|.�Q��ܙXG<O��`�)��3��+`E��f�IQO_�!�& 'D�k�0�
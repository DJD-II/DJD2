    ����          �  ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j����wEj�kB�A~r �x�2��H�"�BДN��á7ڴ �rA7Nm@��):Y�]��/�|��gW�:��Փ]���]�Wd���'��=�a0�a5k��7(��8�t9_����j�sRu�BMM�Dp��{?;b�)�����r/��F������Ό,�]��}��7�I�Ik�H\��Pnd���Y4l?���Y�E���Y�^�c(�w���T�w��>q1��/;� �#'o�Ĭ*�T:�(�^�e��\%Fɯ����[��� ?��`��<�������I̫-��(d:@��C'&é�1D�#)zL�Ԃ�/&F�}
��>o�x��&�ٖ��P| @�$ܕ_�ܘ��r(�n�ٖ�����Δ��O�6*�B��^�,}�Y�U�$eg Z�C�Ys=ܯ+��r��2��T0]2o��i��
�(d�e��J���W���C�lR&��.�Kv6����_�bY�|�� *��d��/���U[��+��p���tsg�3S��*s�c�R
}��}Y�G+ ���Z�S���+�bjN�Y�$W,�����	Ԭ�2��V��{�e3�h���~���#Q�3�Wj�|��H��`�1��u�j:~E�m/g8H����S���Q��(m��%t�H�� ?��������av5�>.:_^�ⳡ��0�^DaCZ�T��R&��B�Lj���j3MU�P���W7��P|��]4>��]��5�|1<G��ͧ"I�|�^|<����0\�}m?��dIg�4�wz a�[1���)Wn�'5�]��n!��h_�K{��U��{�1iLp�զЋ2w�R��0TB�Tm� �����3�ӭb��iBb�,�}�5J�V�'�S�l⃧����!��*ُ!��{���ÿ�[�.�n��˓з�H�k�s��R�H�Eߢ��M�sSP@�G �âi~/SZ�,����?P)0�KO�
���3'����{PΣ�˾�������V�?���L�jsͪ��x`[�c��N�6�� E"�n%a��<킔y�������[���z����J�J�8r�/��c�B�K�%�����N�m�A������P�u1񃱗JQ��Gv���U`�e(u."8��ۚG��7�c�@�92����Cu�7Ը�"��p�Wm����]J�,��W���)ܶD��#�
P�U�a}�{���A(�Ɠ���W�"�U-�z͊n�S�K~W�hM���J�0��]��e���{��"�(��i�M�J�0����㥱m�\=Q���lBT��=�&3�nn9��4�Ud�ms����:�����ǘL�U��ƚ}�Z�P�|~������M0�R���C�A���ߦ�=�f�E��c/X��0���>�s���`�@J��KD��{vi	�ʼp�ӒWȏقd��eIr��B,����6�"leXk(E��.IC�k֭�mi��`�i�Y�;g�LA��h�ۜf�v��늻L0�b��[#퉾��	(dyْ8����"�2л��%���y���W*� 8���QF.��)lr ������n�-���7!T8����7c:a>���oh����Ө@��B��s`6l+�غ)^���#ڏ<
����������f,/�f�D?c��K_|Q&�儔|���H����0���ř�BÎ�'��e�B6DA<9 �p7�X���l���+/��"�y�]:�=@�����w}x�m1i�BMZ���(6�l�
,t?�W���=O]Y�;��uدF���R���N�5��+�W3�r�},ZF����> s���~K]=rk�*���K����ʆ�^w|�����2���-���`�uz��9������x��O,I:$t��n�I鵟޻�0��_�u��)��l{����g��kn��<95�A�=#7#��+��m��@j��$G[8QTB�5ގ����
�B���1��I��j�߀�8�8��2�y��A¸��5�X��	����8 &���F��yT�i"�Vڳ���0�d�H�Gl��e�a�d�W��yͺ\Ղ�Ѹ߮�8r�{Z��cӨo���k�L�J8&�P5�&ݔ�o>ߝ�|�~ڌ�A�m��)a��׵Ke%�����5�]/\�ܐ��x񒖥׼«�hPuq̽�-��7�4F6�����Wg�ߚz���w�N9Y\���������*0�_D�z���ޓ��x�?ɒ�@�m�_2���\>�w����	�L3t���P�M��y[��[@%�uc y�s!�<[�۞��pXN�cHi��=c[6Y��P�þ:=� F��`��th6�Or`�}ʊY*��p;@1��Z�.�ş��z=7M�v;e�����3o�����^y���+oN��`/��O�`�Mƴ���L ��ƾ�{�M���A�$pؔ5�����u8G#C���(��m�s:|x��=[���_��"�c���B����mhW4��K�9�Pk��k�/*r�4�)�͞�r�~/ǰ&J���0�hk���Ak
��G�+��z�������zL�L#��%K�K׼����/Y.�D������`�km_k����e��M&,T?X�+l6� �"��{~�ǰ���8���č��qV�.v���Н��l�c��R�����\>ܼzV��Ȯ���Ɓӗ���#��%��^{n�r��n�2d��q��7"b�I�s��y�M�<Z?���ĔQ�b$s!��ͧ�r,7o۩k������9�ɃT�^��Y��`��7�| 1�����3�V���X�"�]�A�]ŘBV�)��*n׵�5�}����W�l1iЉ\���6<G����hui��P�(1]�A��O�c~xe��۾Gr~y�:-e=��9��[m�%b��Q�:i����+�uKl	�&��@��~`y�~��7K�Y�ĮY*�����p}7
�MV�$�������6uC���������5!擰[)�E�#�9(h�C9{�2�5�W�^�{rf+�w�M�5��B�o��!�e�ފ�B�暻�J�h���}ð����G=Cv�U�E"�|�xC8;�^%hXA���G/���W�3�6����0�(��U	�+or�צ�T`'_��:�	U���@#����+B�hk�c�9���	\�͠ɬmP/b�s.t���	�vlr<-��椺�)���L4��A%�Eo(݈�1�QI'Z��κ1�� 1vC�E��f�6 �F�
Ӿ�ax9��w��ꉃ��սr�,M~|Y�h�9�g���z�/��:��m�y�����Af�-B��l���e����������b�-ҧ';U��5���YAn:1N�H��|zE��#1����Sk<�@�w��`�]V��:z-�Cof��`�jטe�{�=������?��?x��ymk�x$t ���c�n���n�n����\}څ�� 4��������Z	�f��K�����m̋�{c�&���b:�|E��-C��Ͷ&f�).�]��]�/��R�e�^_����OԄx��J�ںA���C؟ό�D�ݑSf1R�s*�0�g�l_J��-���a�8C [H���9=|G�:�+Z-�z���O���r"��k�'���M��@G|���sx"H�bБ:6-n�����6}$%~o�!н�Y���X+[���7R%�W@������!��lȕ�NxtD�u
U�W�AF�q�vvb%���> "�i��<�B[�A>i�'���gTK����*�#u�Y>�lV����0�/饗	�9�㚞y��qb�e���*�uT�nw�ƛbc���C`�0�F�O�+�Px�B��OJn�>���,x����
m"#��p>C���:�?�����)5�s���}�w���4�Xs���!�-%����x�3�K��d��r2[��g�kP�g<���D�8�_��Q+%�K�1>bG<�K@�nB�ơߜ�\�ƻ�K�P�]�/�&��s�W��q���x����w ��>����1�&r/C��7}%]э��nO���G�}-�-��ԫ��V0��3q������P�����`E�����'�-H|���n�I�M3��n�Fq4�y�o"�ǎ/���nf�d���>�"�ʓi}gZ�EQ����R]<���L˯���G����1��+т��r���i$Y�����*h;���$?R㸍�E��.Qq��o�h�tm��h�u�Ke��T������Y*�����F7詥�L��+?�����a�v�w�,�l�bϒ�3�,e
h�S	y�&�������0��5� 9|����	��U%�o]��V/9]�Թl?3���k��c	}g�CH��b\�j6`�L}�w�%�Ʋu��� ��Ή�c�Q!�vf�G8s"Y�/K�J:1�\o�{w��F`&�	'g�_ ��BJ��!A��� �*B�r�4p �m��S�됣�J6D�[��3���p����P:��v3��N��It��_;β�v&8��ǆ��f�m������֝7���jZ9ݿN�|�gb3�v���^	p0�t�ݳm�?g����kO�]��ހ���R�#5�=j~f9�+57�=<��L�G�<�l��S��F*�؄��к��)l�������G�r�OX-&�ȋ�;Y�����{�Z��Aƞ��>�����U��3{J�N���c�*\�q�!~�@0���t-�JF�rܺZ̶���fͲ��?��f�֑���BUX8�YSϵY>��Tf�j�������zl����s[�T��-K(f�]�p���	�$�f_�$nbfk�1�}��x�^[tj���8����A2��N�Q8�:�/m�$�l��T x*�]���zQ[f9�	Br�^N�hp��ܦ�ēe������~"�muHήܵ^���
m���,��(t�u�?�3���[dȶ�b����2B�0?�Ow�F��!3����	^�H�29>��~c,���F�p��Z �2���GG��ov���~��6���5!���0w��eO�?�V8�B�y�l��ȊA]�	��ٲ�{�q��H�H�����NA�#53�4�0����i@y �ӝr�@�������0+�I��p���2��\����<��Y� 
�x��Bg�/\�w۶���?W!Kq�_{+<_�9{��f�7���k���|���,H<��WP?����v���޷�ͷ�=���$N;@��P^�/vJ53�Q6���%�����>� W|��!B٪Jwr5�2�+|4��̼O���Ca�����M�E�H�0B�d�zAc���.��Zȣr9x�a�`�i�u�v׌�My��n.��/��/�c���c'ak��UC�{�#^l�*�[�����'x���^~��ցnoa �0�yq�
E���Bk�b�)�F�g�����;�~؂#�hĽ7F��N��6�x I�J�A���)��0�����p�Y���=�	Z���im�k��g�'��aq&~�iw� Bbm8��3+�\,�n�IᇛA5w��5��O���RH��ɗ�;^QB��<��a��%��H��YhT��Ϛ5+3�;�I�_��>16���H �*h�^�u�
�t�,|��p�(>M#���(so%��7�rc��9|��F�������6�T ��,�N�{��	�Xʉ#71sm��{vyD��Y�^�S���7˵Ք\.���H-�:��J��V�Do7��
�"v�m��W)ӵf�x3i)�Fq}��W�5D��R��j'��nA,쾚1�B��w��uu���B]?���`���Hv�1U��{Kne�IM��fN�F",:5��[2۲=��4���������0Hg
^����@&/a�����6����1��S�hh��a6
�k�+�>���*	I�����cBd��*{�|l/�94	�xl��NF?�sd����a�9��'�8�o�E���W�6��+��׭�\w��;~��4w��s�挌�IyC��o5���Ύt�ive���e�4�х2�gaFD��'�-H0�HMИO}����#���LD���n]�*q6�*�0;�e �V���l��G�{%iQ�D�Kd;�~*��-���;D荩Y���[먠6v�_SAaB	@sRݝ�	�fF���N��{���9u���-"��N�t9Km<6б~�����P%��@�߹�g�.�U����v�p���빑�҃U�$-�坨m�~�^s� �"�y��X�5&��_\p$J�%����;Tb;��ph�"f�b�0�ľ'o��P6��E��v��7�]����8�@(Y#`�����*{��~Paü��%�<������<9��N4W�V��K�B�Q�1�v�eY�4r�����kB��Y(K��1F� �{6�*��@����#Q��g�H�����9��Nȍ��Ƚt�s��"��G��y�#��Y�(y�Wbë�L���:��Q)Vv��h?�����
�7$��Hʚ�ц=}��:�e�*HL�N���MY�',| X�C�ě����=�?�-{�[6�a��:}�%5R�^g�ZE)ƴscto��'����V�:�vj�S���p���t�̳֊>dw{�����G�'4c���S6���u5�>&��;~� �>rn��χ5P9~=�@�i�i��ީ5����o��k�e���JDo�ƌ�)�b�/!���X�$��TF6�Y`g�T�醜����TB�Zq��N�qb�a���8Cu e>��A:�1���}� .aG�G��z��'�|=)T�8�����C�}�(�^��|�p�&jBf+]*XOM���v]�~������.��&u|ăaZ&���p6���Թ�i�߼@���MQ� ;Zc 8ُ\����ީ�א�'T�q��׊�@�3�Lc�	�j4Yӗ���m��r��W���t^��x��]�vn�-��!v4KY�r�A2 �ƛ�i9eQԈ�F���h&�Mw���J5ķ\త-��2l������ �"��I��V��>�F~�ra��?ObX��*߭sԨ�
3�^]���8�PX�k���k�o/���p���ށ{�8��Bw���1N��-�6���:�h�<)���&�?b['��]����Aw��Hc����3+;I~c쬿\�V�L�(g7z���CF#�͓k/���[��׈�̅��n��n`շY57�ot�:?�樳����i-��w}�v�n���5qr]���c��a��h��Jn����)�?�|��1��/Y��L$�̀%���p�wX;��؄���9��xQd�Gs�z)�I�b�٢�2�9��m�>G� �V����H��#{ன�C�M�G��ϱ��{�5�ȋu���3��5��2������;�Y�z��6���-n�<���� 
�C@S�6�<'���ee��t�Xo�������{!i��ː��+���Hl�q98C�Q�.$6��M��N�JPL��V��{&��icR�(H���4�'�S��x2�/֟�|�:
U�k�;�x}���:nNg���o����H���M�9㛊�����/�%��U�S��z=��ř5v���)��}J�QG��^�%���Ve��T��,��V�݌=S���]F���#�.��k����y\����w|jGz�$яr�����XT��BV	������� �>����&DؘQ!��?�R��]ZAS~���,7(�*�~D��$g�8���3��ͮ�	��w����<�P�2Y`����C�Pi�I_Yq?�R��k�z@����5W�ؔ]?����_՛�p����$��-���i�u���wQ�*���_�������7�$ƽ��9��@��-^��
    ����          �  ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j����wEj�kB�A~r �x�2��H�"�BДN��á7ڴ �rA7Nm@��):Y�]��/�|��gW�:��Փ]���]�Wd���'��=�a0�a5k��7(��8�t9_����j�sRu�BMM�Dp��{?;b�)�����r/��F������Ό,�]��}��7�I�Ik�H\��Pnd���Y4l?���Y�E���Y�^�c(�w���T�w��>q1��/;� �#'o�Ĭ*�T:�(�^�e��\%Fɯ����[��� ?��`��<�������I̫-��(d:@��C'&é�1D�#)zL�Ԃ�/&F�}
��>o�x������z���� u�n��y����q��R0�y��%M<c$)@޿P�u�\����%f��s-'7��M�*�6��\]�Xf:����*��W!�@�
v�\�>���8��1��O�~�ٲ)���!�y��gS��Κ��~�ۼ�3r����8QL��h�΀��9��S��r��O�0��1���i�d|��$hZ4�N��X�tǌt�0Y����� X��RrE�"�s2'!8�ă��z3�{�A�Q�ql1#:�T�Gm���'� iBV���/Ή�E}H�D;綢Y'��A���ڴޝ-��Ov��v$���1�B���
[Kt?{�����:nո�:�T9]�7UZ�`D�>n�P&"���
ks^�=�ӓ����{L���=�ȉ��ˁ%������G�-��f�"U��5Ȥp�nv�PňH��po�D�`jJ%���"I}������ mc7̰��δ��އ� N��lH%��cл���+6�Vn�Y�(�Gm�d}���b��k���3�B4p�_���ډ�y�|730ʿ�]�EQ�0ܶq����S���~g�{H|+	Dl�,�D��e�[0� \}kʆ����+��ڼ��RT9u�J�!�i],ݗL���w��Ol]�$���Ôs��+�_� z�'?++#�S�T� ����BS��l#JH�5n�y��П��΄��^��-��'���D+�ý����v���aH�-���V�ᢶ�φ�s9���4ǦL�mN�՚�ĸ�o�X�m�6Uӡ��KB�����-V��[��)c�x�X�+=��񴗜$�Z�T�,,;� ���oǑ�C��4�ѫA�xBjKE���0��?�W �	vi��! 6A�
�z����I���U������������ӫy$���'j�K���]�1M�|�I)Y�8�Ϝ,���X,S �ጎ۶z	v��_���;�F
V'�5h��%�;���:��C����͞��#�Q�.�2�sW���^�8�O�s�$�U9�x�'6��ﺩWwib8�e��v�z�g�tz4<�l�
�ɟ��uk����D�vm*'�{fw-&�X|���X$�M��n�����*�W����k[��Fn-��=4��P��]���1�x��+����P)I��4-'�@�ϝ�\�}����4�[J	щ�uxI�H�6��?Vd�U#���̭jHd�7���N�a��^�kmC�jD"G�h>��D
\���؃��0�3���̳�z�ආ���7R�J��!��,~��
1�Sm�ɸ�C�w�v?�i��� V�1t�o�2�]Pg���
��>6�f}j�� ��M�\�H��7�J0U�q�	9
�H}�rЕ�{�lyřQ%Pt�.�U����Q��.&!��v��[��	�!YV��PfV}M�������Y1Q�BT_p�v�p􌛱	�)A��MM9���)H��9�ԂW���:&r�١�V�y�e�(2|��@dX�ʈ�>�Co+��ԓ�˘toY\E��2g6�	���2HǵWOR�c�,pS	^&�V��A����6~�p����W� +���e��P�z��|�C��=�&ݻGR���k��I	���� ��T.�Փ;�/Y���	T�g�~��'�%�Ґ�� �3�,.�]�R��^��7�{�if�������sT��[��<����)c��D�y���-�k�f4�|�e�wx���sD��_4��ձI��v��(�ѷ�f�L�D�h#��X�G������.�v�ż�L����,A��n��r`���j��)z�J ��r_c�{��D�kd�7.��!��������-l�e��[F]�H�h��B �q|�Y�AD�A��ߖx��Z��QOd�P���./=A����[�(��GL!��'~l��A�]���ڐ�<-��;�m�sg��53�*��⣈Nʹ��Ɯ�!On�!��ˎ�r�R����{�L�Vq��'�b�z����H��Q��T)	V��D��Y�'����|m�Pvs) �u�3ʝ:b�^Y��@�6m�xʈ��5�C������*/��_�Ĩ���,/���d��Ͳ�14��
.�~Q�}��u�S3;p�4��QX`�b�VJ!mT]ф�K%���Ǹ����3��~y�]���;�fE¬ͯx�B���Q���]� ���Yu?}Ӕ1��t�&�n�rݝo���GwK>Dd���S��Wt���XG��^�>�˪�D�N떲Hi�ڈ�qp�� �Jng��%�G;9�jƝn��L\�T��ϰ�G�M��Ǳ�eT2�'��=ojR?0����x��jr�<o�����k �ȵ�����+��2�"��.�_l�R=�%s�����^�"�\���H-���l�).S��5�O_)^��o ���lcŹ�`���R��f�hnS�XS� p�����I�Um'/��Z�:R��xG=���;Ā�+	j�J��:R�FjxDr�1�jm��*�P��f]=�At�8E�=�`����-����mVLn��N�,�/�Z;��1v)�`���&���J��d�!<h���YA��&G�(]�9U0�ț��u:oː,7�?"L��%�K��������C����) [����*z�G�Y*��(�1U��դ�3VE�C��~wr�+)�C	7jgBAC�9&[4�f����Q\J�#\H�N�A���7Q��jm̫h��m8˰�;z�)@�}�O��~�A4.�3X'�����|E`�]��X��+dURGt(��M��+;տ�.�V ���-��Yć�������0�\׬FS4��B �H�ȤRp}�6f��;uI�KB�^�F-�Κ��rF���g���>���������dQ���`�����k7$��;pR�O���,[<�RKQ�0wgM(ff��^>� i/�����j�:[���E����N4�?�Pkڜ�Kx���4&kUf���r��T��"PJ�B�ó��n��yB�p=P�f��qL�#�#m����;i�%*�m;��ע.�	�r����2�oFȂ9�f*r1�$��$��.:�o ���b� d��dɫ���.��T�ܪTv3��T����#�%��Y{`����Jb~��螳<��^0��`��^��r��<g)�M�����
�N8�y���psC�S���g�כ��� �W9�P]h�ӎ�������D�?58r�J�C:���{%!�Q'�ȷ�B�[)#�~_��93��U0n�e�u.���p2�gH�s����x#��H��
4!�4��}D;��D�,�]����hlم{ѻO�H��Ff-�b �5�a8o����n�w�Q�6�����8T����?7�q/EA�5�ޭ�Q�Xxg��YTH
�����QCzMa�Q���mH��M�`���)5�ܹ);��]�v�Q�V��<ݛ�N�r@��sN��MT��a���4j�7C`�@��>�w.c%�Q͋�xJu�D�q"Ē��@�TlF_l�﫥J0O�f�J�+�����NB�U���2u�-"u�A�,�|���6|�ܫp���gu�0�<��ܦ���ǔ��>�+p�BZ��::�9gL�w48:m��K_?&@�Fi�}R_L��_I9���	R�X	����V��~*��@��D?i�6�CA�A��ބqY�Ls����Gy$�N绎��#֣�k��.w6��D��5;�����J��&-m���$]DY%D���z��|қ�U�	�%N`����:�J�7u`	����7�yE�r�v��I�2�������J�R[�p&�|�
��^ڷ�	���'��(H��tB?���!���g�M����U:Kb���t�"�eܓ�;מd�&�F/p7�;��e��3�Ex�v�'!�6X8�`܇���b�6����j�Ӻ>n�+�Ǧ'�[9�{�_��u���-N8�5:�ʮ�L]~�^f �]����m��}KWP<aiϥ4��x<>���gl��Z���j[�]��֭Z�4�́�&��i�s'��=/@3�X�2�,t�(7��:��q<��~҃o|����)�ww�D��Pi�C����mC�n��RQu�P�X-�*^��>aB!J}��i��`�~���Fr�Πm�^{�M���NԔ�oXPlH�g��p�"�=-:�͠��~�?���\�&^��xg���w�ޱ��"�}]�e��Z.MV���'�݅��~��M�(;�`�OW��s]w˹�rZ�ڛ����P�{��_h�7�_���W�7�X����g7�$�< t/�W$��V��_���,��9}~dڢ�1�C_	鏚�Cjhc�yn���s����B��{��}�Y�}����-{+��uo�&��n)�m����/��ۉ0�a�i
MY�Ȟ�Α��4�a/��WRÞ�I�È1�2����t����O�L�Y�TPm_���?��WA�e/���>Y�W�o力�Y�p�n�|��H|>0k�&^�'��|��bs���F�]#���.z�޶�2���M{��Xʡ�_����pk�V:ӑp��换ÑB�� k���}O��۫eF
=��Ԝ�t�2^2tY�IuA�]�T#�:	�sh��Q��B����%,���� ��%�.��|%�\$����扟����~o�/������]ÑLፑ�E��.�J)oc����dH�Oɝ:6*����s�"�U[7��|���Yt�[��C�+���HM(}���,̊����9+z�I���XFG� ͱ��*����s=���	�u���
� ����A���Hbҷ�#M�T�Τs�F�]��z�R�X�&��TPf��$|ҽ[`���`���{׼wn��5���s��y�NM���鱂�͈}��q4�i"��� y��w��q#�p�(�������@��p�jI�N@���u3\$[�6�湼��8Դ��ƿ�{oDīnI �
I�Bxr$��ҟ�Q�Ԏ��Am�]X�P �-��x�.q42��O�ݾ�'9��O���
��vc�+ͩ�Ʈ?hiiƮU���`܂z\��_��q.g���s?	�57��C{���7�l�2Y~]�O�~���S��5�\'..��d�>0&�uLXRf��{�_��=w#����rDnȒ��q����)�A��c@;�Z��ֵ��ɓ��+k��e������Z{�ι��xZ����3宆�l���i���u
6��/F��x�� `�9v�-+I��q��I�2Y���m��mӰ��c܄�?~��O�l�K= y�e#�?���ѕ罅���['9H�#�"���q|2��)B��񾸼���_l\n�@��AZe�{�y1D���a�A�����a���5"N���n�JV�d�A��ә��w��0����L��u7\,�"cOW������,�f?fSu#�yik���A5m��B�ϊÒR���W��1F'������ث*��ҨAO� [�rʓ��"-e	��[�����:(��04:,�������a� ϻ�X��,�M��){� ���6|;-���j��}H�v^]p�&�;}�ދ�9�l�8{��8�빞X�ݔ��B�`���^���<X��q�P\ه��&VUM��,�T�P�nk��О�h�e�}��VQw"g�5�Md���k�E?��Awb� �y�V���]�X s��3�����BP�#�KGEe9�+�rxA=O����tx�'|m�4��0]87�F��1�����M�gDQ��K(뙨b����H�A�D��+:���b����}�ⶏ0�ۅ�\\�&�\Z�%��_�2���u���{���';�Ӽ�����H�aL/�眉�@���y@d��i��0R�)VV�C�L�������x��yq�%�ƟS���ijM��M� �ٕ�{��5<j����_��hU5U�C)}l�c�8YT%�cH�`�	��\F!���	?|Nc��)̏n: �v1g�Q!�_��U�Q�Y������$��hi�Ư�#�!��V�~:�m`��� ��?�jo�H�gl�{�� �*�������K� _E���=-m�o�g�x�����=�
�NB�O^��eλ"��>�T��膧���s���A��'���[�u��x�W���)a
������a���%���\/6+��MER�����:j�^i���|�&��FsO��;-�y]tׯ�Ʀ}��A�>0^x��B�%���^���5�W��������ʯ�N�WEZc��X�¼�V��%q'�I�E��MD$f%��~W]F���h���܎e�ޥ;�[c�&]�]���d�t`b�Ͽ|l���n���ނ8 `E���gy���QIeq�*���
@�Z��ω��5:ߤY��Q��l��á,��Xr��̱��:j:�H��
o�;K�1,@��x�p���$�p3Cy7�&�.Σ$}��_��]���rme�|<Ƭc�;�Dt�䮉��F���Z#+���CU[�3��[fБ���}7��>v����&(����(�̏�	�D��2�v����*X&U�y���L�*H	�/d�9��%�'���P<8P@^�����^6��6��G��0n��@���Ϡ�U�!ɋ���w�e�ߜ�eK��u���%c��3vˢ��&�t�n1��� d�� �0B^z]���)y#�@�⿌���cA�KҌEĔ>���bD{�=m�E��on#�7�
�Y?;#�@wך�k��Z{� �hi���.�u��f�U�АR�7�W�o{�̻������p�W{������ +	��C\ݬ��%����`��$4��4�O\r�K����7,L�:Z����L�^�i��`}O��}�C7�b0Ҳ籢��GC�,&��T���/�9���H�����un�Ѹ���9,O�u��������� ��,Ĳ��FѬ��B���G��ʑ1�*�� `��!^�
��Y��|j�:�Xo��q�<�H^|���:�= ���C���gu ��s?)G
z�~uA���$Z�L���D!�����F��Z��m���&��5u`B3B��`4��ب��B��z!��ܮOv�'B�^x�%���*��!B��D�5>�L���C}^�����d�ω����z!�|��O��W�`�^}�cw���Td.�W�Ա]�ۄ['��z���,�l�\�}��d;}c�M��n[���;E�ٛ�$���d'y�=QO�	��/��0oGh���G'��`�$�q6�l7hD �>'�ߋw����H��5J�I�!�6�-�g
*D�0L]}Nֵ��/T� �0�S�Q]t���Q��@<��$Amo��tI�gP���Ft�/��]I���>y����m�u	��F���*�(f��*��x<�؈K�v�e�D��JN�VjB�r��W�"��k\�7��T�v��׬Z�<sO� Y�8��2����klN��l}%Nd	�5�J��c9Ҋ���@U�W]+q�ܰ�
    ����          �  ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j����wEj�kB�A~r �x�2��H�"�BДN��á7ڴ �rA7Nm@��):Y�]��/�|��gW�:��Փ]���]�Wd���'��=�a0�a5k��7(��8�t9_����j�sRu�BMM�Dp��{?;b�)�����r/��F������Ό,�]��}��7�I�Ik�H\��Pnd���Y4l?���Y�E���Y�^�c(�w���T�w��>q1��/;� �#'o�Ĭ*�T:�(�^�e��\%Fɯ����[��� ?��`��<�������I̫-��(d:@��C'&é�1D�#)zL�Ԃ�/&F�}
��>o�x�ېy뻑Fi������������_�\����*������~��?~�Hޱ"�yXZC������c��28ג��[�u2W�h�C�bN���*��m��e�%j�k}�"��ȆAK���Si��G#[���>ur�UԠgCF~L���;�i�yqj��^�j�%;�o�hg�#���pn��rË�'#M�^ݘq��fU��|���Q�h�����.~o7��m%��⸞.Z��_�r�����ά���s�sC�������/�6�۩�݅����6�Gl��y5�^a?��-s�(e��f`|����p���3��E�\J�};�ax�����aw��9S?�6��>���2�e�`�C�a�VL���S���5
�GpԂ�eH8*��9�Bʤ�WN��9A�q�u�ɇ:?F&�6G@	�M Ѿ�:�-����]z��̆��%���p��Ѝ�K��{�=���ۻ�2�ҹ�2��h]3$�6��6`�5�Y?U�
�K�ճ�%5���#uk�)��ՄU}��X%���D�y�S��c������H��{D��jl��l��¼�3�7e��
������GUm,��͞O���<�hS��o]��s@�~�ݒ���AR�r��B�'3h"�+ϠFƴ.�bkm�.J�P���\��!�Pw�l��gtM�L��I+�~ɚ5y!~xͥS<[$�l��TW:��'�	S�ÖN��k)�+=���'l�vZ��
h�3��ȿ~�9:�z?[h�ה�xl8�V�QCK⋑�"�z��M�9 �M1jm�}_����2���!�_:����{EF��Af��J3)�{�W�+�c�м����f��O��vJ�$��P�א�]�m�ZR]5 ���8.����*������o��&��ݨ���x�dB��u�}D��?tugcq�)��F�H?OF�
����(L�#�]Fb�� �2��J�ަ�A�i���u
u�uVX�0n̿�W��-��8�́�ݪ�+���)��Cx��vd5TD"B�@�b�ā�{�&G�Js�1HG���TGp5�x.岶o�>��o��*t�`j41�c���hw&ʝ�C�P������;
�+��=�5�.�� 
��d�@���A�)���1��U��w�!T�ς�x>�����/�� �x�N6J3�ÓY����`eo�i7�P�A%��& ��r~ړ��A�@zJA�z�k�rB���9ɧC:zḰ�l:ЕD���aJ2=gE����W���'M�BȠ��H2��!T��P�bڐT��}�8����#Avj?*y�2��=@�T~q8��\��h�윱@���T�M���;ů�m{�v���b)�b�Cf��O.?�Wݲk[y,�2��Iq��\��vM�(� g�1�Y��[�'*���5
��VS��Ȑ�Y��83�jY�a����H�{�ك1=�ڟf�˳�ݻ���G$�B�m�J�N9Q���&w	s=W�$�T�`�m������q��[۠_T�R���č���]X�p�o^�5��3�8��0�[j�wg8Z����������Ş�P���i����}
����\����.''9�]��rĀ1�N��n$���L���;�F��4��B�� 2 �vV5&�* ��N����6K2���^����Yw��&z��JPy��/ƭ�Iy7��OtG�Y�H��~k��b�p3�:)�싗�h��� ھ]���n���+^�>�ȃO�M?s�Q��*�h&�q_�Xq)���r����c�a�wK��΍`)H��Y#�7�We�zWR&١�a��-x��q���S����v�g~�;}�� ;� ��	nsoJ���6.�k�{�Q\P���)�]��}O�z��k�ʇ�2WD[��<TKp���מ��֘P�dr���4曻9�p�&�L`t༘�ez.V_����mK��:~N%��pL��X�iq�\���ya������3���LA����(*�@�}��5�Y����� Cre�L)ū��VEcT�o}T�̝�̃C����ڍ�h!������t���J�Om&��.���-����¸;�]����wL2������G�kF`/�ɂ�_2�j�'�~�d�#� 5Sj�MZ�:�z��9�mN-b��O4�Jk�T�d���V��[ˋV,md�C��ڗ�f�1K��h�n�:���^�T�(��o�4�z��qx/(�B-5��2�x�JK�[p�!�����Ǉ�Һ\����y�8}���Ô����y��L����㐪ß��J� cߌf��)>���[���znQj���"�"�߷�/n�w�z��3)��A�u�d���i�#U�̤�̐���R�w����!aUt��a�Ϫ`�s���o�9������}�\*�:�P7 ������Ӊo�^���%*��)��π{����E��|@���R#1���H�./VHh0�ja�w_H>�֠h9Uv`=.�?�!�8����!u,����|��V�����;��d�������K_�l����FP��;���cs����Pk��Ԕ�|�ݳ��{�P�`�%=�����)��+���	9L�B�Zl�����b���7�X/��p]�NVU�,���a�������#RI*z�M&lMs���̅I��P�}+с8���{�^!�,k�A�H���X~g-�ϐ��Q�o�f�6�ؖ]��O�.G�*�Щ�L�� 4�R�	��[e�.�F�S�,Th�8�X�N7�H��>�ҍCW���}E�ʑv��&=I��b���,E	,qYRl&C<����+�f�ɝ{�ˡa��EB܁����xKƮ��@+{��;Q�S����4a�I�<�����I�]u�BNӠ���9GJJn>��f6d��� ����C���e|�e'(�`J����Cȗ�:6��<w�隯�]��4�D�2����{E����Z�Z��e��� ��亮���T�h-Û�5�f'*�!�0�.#�q���("`��
ω�0�*�"��|O��i�<ise�8*��"ב,˟T�@�A��%�3���O뻔��-��zBi����b�L���)S�f�)��ig�aO��z��9�����gS���Ē��쀭�Gi����*��L��Er�pd̆�nя6ҷA{ש�ܦ$�2���q%��Ё�X������J8C�^�M��o���u�?�v����ڇ{��5��h�%f�5��)��3U���{%�O���YXz3>��ȡ�u�~��v=}N��o�S�f�����$��͜XUfgU�a�9��$Z�T� oʣ�Rn7���VrM�P�XIA���v��>�:����������Iv"@�>Ihn.�9����i�ʑ>|a}@��ޝF�c"=L�M��Z
 3}A�%#g���
��N�Tqs��@m�Fp�\�|�,��Lo��}��r���B�=YN�>��#���L��	2�]�;�%	j�T�T��:�NƗ(���0�}�4ջ�mO�\��B��p;feH�I?q��F�7����aq��7��GR�aΜ�D��C:�����v�FGi@ej�E��:�ki��ڥ�{9�p6�� 
y?
����0�axP�6o(AI�m��,P��.(t26}V��]�=Zc�fwO̭.2��{�� �oRn���&VǕW5ϓ"N���z�{�.�+�.@k�x�b��w\r���7�P͑{H�A�����>j	v�7\�������H�),؜w���`@���5�����H���>�$��a\:�&�3��	�&D� �q�0z̟�����t�i��oBUWys�T!��X�n���Á,p��N@��m%֮��у�ʮtAtP�= [B��[Y�Yj|�;=��y�*�Kc�i�m@�_&{����G��1���7A�4��d�vt�����zd͋7q�wRQ{�:B�z��`et:�%�cÅ.�������2���6en`��A��z�k�H�T����<��С>����Y(�CX�B6��B3&�y��o��eA�f�f�f�u�SV|l�ڋ���y�&nBf���W)ay�Pi/�%��m��ڔiԡ�tiC2�!�U�A�Y�y�I�/����{�*�*����g�2��� 8�l�R�˂������D}o0AD-��_��tѳ�*/����%���2�-�+3�n��x�WpE��E�n�ݗ�]��T��B��c�;_�l��%��ͼ����*��_,DGիwkd�ϡn�~��T�Dֻ�����.d(�/�7X9Xa��!�v�?@'�����'��J�����ZԦ��̽�Sh�7�'��ž����I���AM(uRj���Bg��v������a��~��v��@�)�e�3%������{&�r�?�[:�~��n�J�	�g>N��X@t��w�h�q� �qVM<�L��@�/r=\��Sy��g�s��64IxބZ�g�0��������x��8ۃݴ��M<ӑZ���U5Ʉ������V�"(�`g�}$��J/�*�Ӓ|�5��fi#�5^4sCc�����*�r\G���W��ڙ'����|�	�o>3�g�7R |���F����c��O�8B2��%⚺�dIiA}�M�,_�j(�8��~<.� [��F�h�;�5"3�Q����KH�>@N'����H���f��]�Um?���~�<�.�3QT#i�M��b���	����\�7�;�ܱ ��N۰��(�H��� D��e��] ��5��� O�ow�)��`�z)�<rv��h���Z��x�S��Jv{ !i��Y���>����}������׼jc�)�W�m88Oq�Px��#��bDEÒ�<4���ڍf�t$��5�̾:	����x�ߝ�`ۨM��e�(��9�}�t���"��������\ �H)�<9���\~��zuf��Q/NK���\�1	�cCKx/�~r�/�N|��U�~���.h�-jo��5���� T��s�]��d5�.�F�L��z�!f�9)�ޗq�,.�7���t ��J�Y̚�OvG�w�������4�X0^��Q���nOQ�R��쑼ZV��������eM�B�DQ�'��%�B�ȃvI�th?,�z�Ui%4A�d�a��A��:�7j�d�/sqڕ�{�|R\�ہ����}C:�ordQڙY��)�" 80NP�D3�B;�Y+�I1t hXjf�Q����np�x�*�7�t���uk�5>��yJc �a�R��u�����]�C�ֻ�`�y
U���ZP�~��6�g;Бl�Q$�>qeQ��������	&uc5�=�/���p���|��(���=���]�|RbU�����@�@M�U�ِS��u5������ap6��������Cn���o>CucnVp�<C?�Q�\p�'��uF
yn\ט�4@�:�lj�oLP�g-h*�<��[�{�*��f��C7k��_���t��>�3F�|��j��# �#��z�'�M����d��Ō�I'�����L�pH6�giMn��\JT��h�e�A4��,��x��m�v��П!���ū���� ����|��2�ƞ�a+�������O%��O���%�b����W��(��9�#����q�ߣ�a�
�V����7xI�dI�	ݴ�*~:]�E�-�<��A��%toy��'�\k|:C<���r��鰟�@`���(j�mtNA=�i��C�`����6hv�����p}3`�;g�*z�ȿba��V|�_���Ujs���ɞwqs�`����^�m	�1Yy,�'��� �d�\T�9��l��ga����=�\T�[V[��ۯ6�'�`kćH�ٓ~���`4E�u3k[f��v�:��B�p̽���y�Ĥ�`g�P�Jٝ�>�jBﰞ+G�t�J��2��^�֝���+�����1�ќ$#}L���<�?�ϬH)v�&�=�dq\��2��B���<:�H��ɜŇ����9x����$������؁v��|�X��4�ʄ����/�u�/� �t �K;J�v�V�����o����O�ܺ���މ�E�[��N.�C���¦�o�����gy1��9k��넀ۖ3�H��*9G^	�a�F��ǃ"L=>/Dϵ!2�o*KىnZ5��F��NMi�<��Ro�N�����2�����~4b��VQ*��|
����kT�b=�e|������m U���̀��d�%צ�3�@���F{5�3M�����of}��ؚ������h�r��@��0�"���b[��M��|�F�&W�H�����X.�Q_�݋�R�K��^-*�:������PE|z<�T���N-t���a�GH�Y�q6���0��;-#�b����]��T�˞s4�b�\zߑ�{��W+����Aq�����iR�����;�6��48�"RJ�+�K*�˝��ɶ>�C呱8d�X�Z���T���r+����U/{8��Քg܍X�ւ�'��/$p�&��\>N�!���4�- ҙ� R��J��I���@��м@6�U�J7�U�MяK4jy)m�f����4n�U�����^���v��d���h*`қ{u(g�N��7��@�+<"�w������q1�鬭r���m�a�Gk�+�`hT�z�Y�PY��������)]H`���*L~�΃ܱV�RW���D��,�Nۧ�f�a4P4#9ݚNg�ȱnA�h]"t��C�ji%�Q��Ђ�r
2<��np]Ñ�K��)�������h��_K1�?���>��{|a�]��s��j������y?�s�D�e7�Z�U��k�����ir�J	~/)\��?��+���`+���>I$� �e�M�a�i7�\qx�1��1<������AB�D��X���4�L�(p(��_�92>2�5n
Bkjy�H���[髿Bݓ��?�"��(�5H0	�l���a��+�2��������F�J�8<#_$q��
,���"(�6���ͺL�J�+��;T����=l�x�n�>�o��:ٵH�廅-������I84��Dz�!����<4ʎ�Q�vx����)eq��[O��C9>C��/~n��X��>+}�`�?ξ���(Z��;��~Z������ުt�IJE�֪��"���_=c���S��؅�(�l0@pCŨ�_Ei��$i-�b��`'���6(��:���>n�v�dsZ�ާ�M�ivKq�1�o^]��ŷ�{^��L�je�����U�eWǓ"�D�2������i� �0s�@�TN栋0�����ל�R2x4��<�W&'�9[�jc���H�<��~�5El��X�0/��'�h8��_2������=@�����f4�|l���l";�i|/�ke~��/�S�l-;h�����Y	�*��V�	��).���s�o�+�%CPq�zƞB��Tv= d,�������c��nt�}��@boI���U���=����&|.�(bk+\��	-W>d	*ڐȣ��� דOCĢ����,5T��:g�̏uê�}���-&	��|�N�Wg�`��$d������j�y�V��������|�e������ �B|[��3����0
    ����            ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j�O�_�S��@�< IǕq��=��9WK1c��EK��ԣ����H�D.��	��T�����"O��#�WJe�l�Gxe}������!�Ea��X{�t>X��E�;E[F&����#�AY�����	�=�F�S�K7��i�ַP�;����Z�u��߮���S������P�ގ�D�D3R�3�����d�ր�^iD�zo�Xki��|�X"\g�}2�-����e����ѿ!�H����E{��d�a���H��AQ�����͘$��aC�-_moq��]\n+�����-�) �w�COdn�)���gHh�4�~�{7f�x0��.��G���SX6���Y�^d%<��t[5��sgn��	�o���>cj��9}Ր����f�R�����/^�f�.����Z�K�N����>-�?AäJ�[��9c��_@~&Gp(9��լ9ν|O���5tsަQ���^�$q!�)V:�{.�g�d��Db� �.�͂��4��� ����&r���Pi���V��;�|�
��������6�K�� t�P�TG����e��T��u�m�WO�|��_1k4�LI����,ZT�7E�C�k�s`Њ��u8�w�<n�,#��r���W���I���A���!i�!������T�Y$Rw�ĺ�T��c�mJ��oǽ~��ff�X�Q=vR���=K����k�T�>"|މ4�ܮ�5#�٘�F �00�ݝ�����1���*�m�*.*�*4�O��#[G�w���<��~�zUdM`�	CX����BlZ�i�ez}��=a��:RC�,��������Hh�k�n�<D�[3N�D��#W�EV ��e[mupL�j�;b��yH<����v��a9�������e*`���8��y	o�vΐM]�񳥪�`���^91����b}�8wZ�J�1
�k�q��z<�dtm������Qq�5wT��Q��)�Lң*�h%�4��
�_�e0e��(�U�k��P~":U�g��ag)o�L����m�`���Xt��mr�$��FJ�zUFȽ�ｙ��,�d���\��
N�i��e�����0U�ăX��a������.U��	$�A�[�*��c��RrF�^�p6�Z;��r��~�c�L}�)�8�s���d��ɦ�,`�&�ԪS.\xL���B�Բs��mﭔ�Mz�ʉ4�<�1`⠢k4B�ٹ�#D���n��lWB�|C;x�y��V&Y�
D�r	6l���g0Ss�s�$��<ĉ�z�rb_|���!�`��T�G5i�8Ī<
(+�E�,y%}:����p�Y��u����X
�Ӥ��1vP@P����������Q����q,��T�B-ޮI�)��<h�ǒ��w˒�s��h v�V&ssy����/��,�m��C�M���y��ɞd�Vg6ַj� \�� ��^�����5��N�l��(�q	J�N���i�|�J	�]vc �A�u�.WaX���z!���b1�A��H�-�xҕ6J�ܨ��N��3��qfP��#�_�@��~����)^��+r T�㤧"q��s4��#������Gۄ\��'��� ;����/���d�"�(��1ڸ���f�0�t����F���l������$h�E'�U[�.�J��Θ<���	���x����<rc rE:��CZj^!h�;\p
�9�X�j�~�s\�kR�����������x�e,�{Y*�n󃇯oH,��<B��M��< >JY5�*��3�g�����a��c}x��0��W�V�C�n�C3��|�8Am�*OQ����v���~檏9^Ǭ+0 ,�2��:��G�o��XJ_.�Y,� ��c����\%������^���dL2
�$�+m����69�@�<0�mP�[��!����_U��s�	b���t8�\u���󥐰k���B�<�kZb9����!�eQ
Cg��7�	Zi���0��m�6�޽p���4�s�`����#�p-h�D��/D
Tk����h#>���\�cT]pr�q.VW�H�!�!u�{ћ�{�ߗ�T�n@�#"���E�=Lh@�Pv��v��אY8���"���H:m���0$�����J�Z�UeKr�!�/k:&t�#�C�i�ˎ��7�,2�0~#�om��A����]���Brn�-��3���[�L����n.$Zrsq�7�&�0��8-���ݱ�&B���;v�����{��KX���R����T\�c����!�I���u�<�_GC��.0T5e���39����ãܰ�Ɏ�uR����` ����s>|�euR�`����;F�-_��J:�災Z_k���z�K-�����m3��o��W���T������'	
]��k6Φ+���q�k�n����h���e����t�3��/.wc%Ó�P�q)��O�⸱��DjV�@��.�־�o�{Xia#�������}A����E_���|!M����,E��vx��x��8h��H{�uu"X�hރ�����Җ�і�kp�A��%�@��┸'�z��^S�Ac5���kr�-3	8�S�}p���S+7K���>QGo�����B��230&=H�?%�߀��u9�㒔 n�; +	(t��e�&�0)��P膑Z�$9���%�Ҁtq���ۢ�5����۞��d�8��1#��Wٿ֫�u��HCTڹ�Au�u�`Uz���"��1�@V����.?�'��͓eQ���WJ=���!��ݛ�v[0
�7E�XO6V�����9jΝS���3>�<�yH����5�o`1�RX��>p%H%v���o��{���g\���ފەI qN�&֌W�S�r�k�hz�1�|��Y���,��܊��XA6Ŵ���̖���Itմ�{`��M)���޿;LIq��X�O�U]f�Ҫ�Jk��\�({k�y���(Y���7Tl�A�U��#M-Y-A�in�>J��8��z�%��R��T�<�,k?�rx� cd%����,���d7U�����K�5�� �e.!�<N��F��ܦqS7���z���Gx�8�{jBa�*(n���V9{�6^��������L�P�썓e�ƀn�6BL�[]l&V:�M'U��H�n�@=<�!¬� >�_����R�)�}���.�!q>��n�f9>s�4��D���M�D	 �����ZtI�:����T<�e37V��5.-�j��6���[�iݥ�ܸK]GC%��Ď�GW�R�L?�a���Z0?��·k�&=l�4tr'�ҝ~�"�p�Ԓ�+�F�D.]Ե��^�UENH&�����h�����PdIK蠺��\��Q���ES�@e�=V��vv�_�>� J��t���W��J�1y����1tW��!n��O�2	��:�n��t�yCf�crL�s��a:���gs�
w�SzR�@y��\����-op{p��i U�(MM�+Iw��d������xW	���l]2�C/Pl�MZ�(��l�P%�(�1<;�U��L�ҹ]j-������+��I��9��be�oB)k���r���y6�sr�9�v��؉c�0$�1�@�~[q7��6s�^f��龸z��Β�({��^���8��z�*����� Z��Y��_�&ކԼ5L�?�\���`�J6Y� U��E�4��%�q���3���Kiپz�ui��R�*��EB9�x��������&i�ID��߸����S��E]@�oD�
&�/!L�niu�P�'��a4Bh�ǧ�w�yC*������v����3����虫��}@QR"�W޸����`��<P����i\�GqV��L�o��<0XLC6j�X����]�ŉ���9<M#���L��/�Eؔ2v-d� ���_g�qP�:��S��!%o�y�j|�k�ٳ)
Lv�7�j/�>�ٿ��ܽq1߹�55�7��@b��ljna�TL߳�6���5�r�d�Zl�)��`�������}8�V��2v�J���A����6� 鋔3\+��pV�+�6Z9e9|�r7��G�Oޏ�<	/
~�4��K�	%� ����ו��r���������	KP�+�A��t����u�����-�	�h'�	|]/1�A���n���}�;6��%��v�(�z0���Y@�n�D��҈'�ɒ!�R��T��V/&|�R~!��*߱ĝ�ȼ��U�Xꦯ�_g�Q�'�Xt��L�l����Ҝ�@�D��2u�f뵄E}{Z��0�;*>�-Z��S�HO�t�(�����*���� 	=��)�C�XI�2��+�=pPީ����$h���(�%X���M�0���2������ՌdA�}#��2��21��!��K�u�(.����=n�լ��|A��asE�J_�9.��=z��B;�i���c`x�n�{��Үi*�1�iΈZ��	���T.��iP��<��=���z2� l����O>Oo�����V�	fͤl=�i�IbB%;�K|��`;U�(�t�"%���[5�v�2>�5D��x�����X�S�1%.��&�`1ɪ��?;ap<k�h6`���s?<�%O�Y�'?K�!T�w79��[S�C���il֔
�ׯHr���0�4{3\2�TT���/h��]gz�ě/
X����EI���Ժ�ΙF\6!p4���u�>��\��h�FA��;�(8�:#���>cv����=4:cb��30^�M��>B�4q��Gf%xJ'�O�YL)}�I�.�Z�!���aq�7��lKj�:6���kr��z�x���\y�����QZJ{x���-�@��	�zc����hW _��E,Et=7O@ �_-d)'f�f�G��v��3���@B�L���&j4��#y-6�(z�S��
B�TcA���g�9g�n>��Ÿ���aA>�MoCC?5�0�/�!�="����5AVkpϽL��������˜����LQ���M9�án�t���֫���5�M����o@-1���z��&���x�	z(���F�H�x6�O���נ��_(#N����,ú�ʳJD�I���q73;٤��>y3n���]�j��� :a�C׊�:=Z%9�� G/�	I�9ɌLD cq�� �⌵������P+~�q�x	�
�RN����<�	���J�T�N\�#Q ��¢z4�o���7+\�͗dw�V����?[����LW;v�~�9G�J8})�u���'*�c���"`@�1&Y�H������%c�M�w]��2�J�� ,��� b�CU�Ds�q*��	k�t�uu��V�+B�.������E�4�.1_D�����/%��XfU�$}�y��CHԈ���&��)qW��u8,����ˌ5`9>a�XK�O`�'� _���F�^a!�͐���G��ä��ܿ��-�k��(��>��f�� �x��}�`R�[JO9Jׄ�Q ���s��6.�IF7�"	l��yx�8��c���fz&Et3���dC
�cNEu�e���U����������5�e���0`C+���{�9�.��>���܈W�x[H�ek'H8
:b�ҩ�I�\!+.����3���/s����=V����s�t�4߰��H�#��"���uJEQ��M��m�b㇦"���;�u-���x��gh�H����X;��M�	��8������H�F)���m:c���q=�R�������JqIe?1gZ�P�v[�a��تˠw�I52b8�Y���S_߫z�jil�K������鞇�#�$��C��.�[z�mR)��7E�wR��r�"T�{�0/R���^7�N<c��ωI<�����W�"��9aa���.pv��Ѣ���5�3��_ ���2�+,e�zWJ�2>G��*jl[Qf�b�I�{�݄&�ʉWv4���1)NZ�~lp���-̀���p��="��GI�\�+�u�f�2�?�Un�� 툏�o�ுd�p�tK$�����4��T�-7k90Qh�j��a��̀��n�$ؼ���hS������Z��0k�y�̖�*�W)��{��w����#�l���	y=
%���B�Ό�h��| ��BB��.zζ�C�#ծ�W��^\��}�H}I<��p�Ys��/ur�/����"���0��$:��R;��}�n�½�hX���kG���+-ֵ�� �24d
`�FYJҝ߳h�h�S�z/̟��39�z�� �N�'O�gg�PZy���1��K��BJF.�qph�pܻ�,�1�S�{߱���;��廙���6��M`��GH�0�	F��9���!H��B�}�.��"A�F�4�0t}�|�B�F>k~���5����_Ѓ�rl�ib}�1�'���fK�لDnC���4��Eo�?�t�Y��7|���4;���DF�g��������c�5+ⷓ5���+���EE�D��1/��=/�s�T�-i�M|�Ѕ�)q�{��(y��������=^��w����)}%_���غX� �A�	\/��=u1g�
Hi0�0ˑ�][xF:f�$Ol���B�֗6�#G����K1�<���8{�G�������	�zI3s@�$�c�Ӷ��T����X�Rѫ�C��Z���O<�'xwE�ĉX��?�gߵ�w�{�z�������wo��4<l�&�����pILr�W��~!�:��M�?l�s}澰�ۙ3�]��/��� �U*xFs�N�@{��f�[����M�%>�Xq�	�D(K��^�'���}��*L�n�ݡ~&��<+�P��~����&S3LohJ���+o��m��4v��(�	���o���A�ۢ�|��\� ��F+�ʋ����m;�֨�8=td�3l��F�I^}m���Tg�S�� �H!�����������\SX�ͣ=[�ɩ���]"�{�:a>L�Տ5?�V��Ƕ:�"�~����Da�b��)��`ܸ�9�X���E�J�oD\�f�I�_�v��x�wY��)5dn0��z���OW�w]�`�oG��rd���A-:#�2� n�Okj.�(�c��҅��,�7��*�+�F>5�Ғ|�_�Dv��	AV�����������RKߟ������3#s-~Gե�.�K�OJ9g�ujL�V"��j���R.k�rT�/�����,#JPW�G�wѶjVU]�'8/��&H�����i�¸��C�{����
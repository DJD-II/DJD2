    ����          @  ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j����wEj�kB�A~r �x�2��H�"�BДN��á7ڴ �rA7Nm@��):Y�]��/�|��gW�:��Փ]���]�Wd���'��=�a0�a5k��7(��8�t9_����j�sRu�BMM�Dp��{?;b�)�����r/��F������Ό,�]��}��7�I�Ik�H\��Pnd���Y4l?���Y�E���Y�^�c(�w���T�w��>q1��/;� �#'o�Ĭ*�T:�(�^�e��\%Fɯ����[��� ?��`��<�������I̫-��(d:@��C'&é�1D�#)zL�Ԃ�/&F�}
��>o�x��.����}����mW@�=����	h��EE���դ��H��"ّ�<5It·�9�U�s��T���$�#=�3ۤ��/�ʆ�����`�UO,�ğ������K[�i��C7��A
{�Ƥ��?� K������Ƃ�z�� ���"Q�&��QTa���d�.$6r�+��$c(�)$�����g�H����ޏd� ���y:E���}�O+�Q��X��;NhԹ���tƎh*�88�D���H�.���K���<z
lvmG,e�����7=��5鈮g�C�c;�O�,���=���2� �`��J�9���ȝǫ���Z�Hl�����v�ģՂ�O����lbg��E5E�����e"���P&���g��W��݇��,Jٔ�78�8m����� G�Wt��[^��� W�b#u#z��׈3�g�掵+ӻuQ������_�~��sV�'��� �\e$8#��c����f'iG
��l�����u�e6U��Лw�����9X���l���y�!����+���]��/휠t����:F{I|rX�� G#WP�X|^f/���������ir~vRZS2�����>�_&}�<{���JV��V��{~�:ƫ��t�!�qd�fck��<yh�l����XB|(�q����糛 ��[@��M��� [�':0i(ť�X�o�Q����Q��2P3�\����s�i-@5�9
,]�IrP,����W�����>�T�h�v�CK�L�o?U�����A�P���A�O&����s4�l��W�!� ��b-�ث�����B�T@��yB�ze8)ne��zF҉�M!�E!�<"�{��J4�FCm1�k��`U& ×4!^~�ળb�&�-b���*ʢ$N�k:���u��[�K��6C}}�����y˦�ֺ[�F)��$��1Gn�åα��T(^pT��b52�3������S�����@����'X/�<�:x�k2�D�z�k�'��\̥R��(��ZS]���ں��p�Vxc�U=�~U8<0�k�pF����Ո��/�q�lo��=[%2��V^���0��:d�	Ȇ+%�/�j������,2�w�@�!v��ϫ���5����������p�������J�*��N�H�CZ��TUR/�%�`Rp/���I�J�|\���*�4Ϧ�=\(���>{3`ѼpuAZ��3��T��E:2�4l�wwP�����I@�1S����b��V�y�2��G|~�w�9I��:����eY�巺S^�w�>[��>q��啝o$J��3�4��I��C�if'r
�u�I5��<�7�hL�I
�i�6�1j�~���R8��86MΎ/��M���z�\f�2�zN���S�1@��1$/R�5l���J����W4I�������1����eL5/���l�%Ԁ�Y��èS��U��hG���%Do�
�ߑ��h�Iʆ�C�61Fg�31M=��t��M��7C*�sN%��1�t�{J]�̓�˅��M� ժ����mi}3b+1ϵ��[-l2�@�YU�@|p��M� [Pi�����xP$�����WO<�%jg���HV��F�C��Lc5ׁkc['��ߠՍqu�Ա��38��0�*�ܒ�y%h���I<5�c�O����ހ����+>\�k\��P�1hs>'��0h�)	���[[5K�0�m��ٍ�!�4�Jf�d�;u�d6~�����0N�@X�3��\'���"G�6KL��s����Ѿ4&n�K�o��h*lY�e (�� ŭR��hD�f�a�l�����h��?l���A͵�{áF좰j��Gk� `0���!�V�H8q�_qL��E����)��¾��&=�O������?��vTa$ʧuFr��������������&^ �؞=$�+#���[W���$e��煥D��t�
�<��܈�����4��B=l�&�ڋ��z��'oY�����\���tmι˥T�8�M�at5���jc�YH�~.���A=wS�=P��^dGk��s3X-09��O~jT����y¹7�t�F�>�]���~��뫨y}��<�X�����S꤬��ZV.���o���h�P<�|���_B��L�܂�GS]�K��ה-���:��W�=���eȝ$�/�Ceu���u�`�6N�
��%?�/C���g�]i|*�ΈS)��y��I��������%��˝��wS��ZA���0�lA8�0׏kKr0�Ѣ�5���l5O��IX^���t'�V��o=t[�Ew8�؏�@�LصO���Z}^��L���Bxqȍ����q��s�������!%�}��X0 �6��!��C�IQ����N�k���71��Q؅�@Hm:@U�I�s)��a~ͧ�m�.;��TG�����`�ɫ�/��^�#�YhF@C�s�E��W 7}����<|�	���Ɵ Ϥn��&6��g��I�rS+���j+F��h�����,W��M���ό��*�`��b�ꆧw�,q+� i���+��|[��f��P���Uj5���B���13lnaE@�Xϔ\��U��k�b������0��!�<���,Ui����6�%FR�3|�ʽ�:�+|���ѷ[?+:���j^bv��<�)朰�����P*�=��5J�E!<ڈ���I�c �*T���ܭ4&�oe�S��'��#�$�Ӛ4Ep֨����Q[<[�4���!^����|n~h]��n���y�W�X���W��	s$�6X (U��>����)՟�rZ�jRc��B�k�0�N�O��5�m��sK=׾A��d7(j�9������	qAUT��z��x�I\p�aqf�	�y����ϣ�;�ؑ`������S�P�NKJ@���5����C�O�jv��78����pF=x�eJ K$��׼�T|�[_ FHMWʀ��r �w��B"�$2B>E�SHL��#n��,re������`��눯�rQ��I��-��<�O���l�0u��1cQu�
��,��a����J�l�e���B���,����}K���C�b��x��F�U$��i�fr�;�P}��+c�؜����_ ��@������"��o���D�ӵ,	��4�{������E��	dz}ƾKBغbj���KL���3���ß����O�x?�V;�kh��>f��}�33ۑ�=N��7ɿ�l^>�0��c�y�P�[�U��-��j�Z��
Ĝ��nɳ��]hx�A�aj�ɟ2a���7sm���K�gSsV��ڪ�]h��^�M��~,M'�u��4��/�5��yZ�w�_ݺ����k�b涸������:o��+����]�1J	��#X ٢�By�2���I��b���iK?b/���v��lB�v�
\���v�>�u�1g�p�2 �g�� _k��i��9����v	�GG_kD]M>O��G����^6w�?�E��_�o��{����ډ���f�),>�ɸ�:��|��t��P���U���X�?*���$���O	F;�f}�B��V=��1.��U�@�dV�h\�ψ��e���;��`� Jah1!�[���5�Ķxg��B���s4�v��������d����W��"p�Y���^kq�c��C�����l,F:�f:3〒��`�:\���G��������j�@ה�ȱ��%T�s�����:4���=`�%dp1/�7�^��f�
6[_�'݌Y�[mfN�xs�J\��54��){b1(�+Fs�U&���F>�1�����	&���!*ӛ&DZ�������w����|�UF�hc�R�`e z#�g�T@�@�h3d\ِ��8�[�ܵE1�3ڡ{����ח�J�z6(����I>%D��+���cZ�)r��V�n�	a1�N��e������&����TF�>W����o�XG��i��#)�#��Ê�'R��cQ���9.��;&���7�|5!�œ����f ~L�1g�&u��3�݇;"N��?��7��,���فyk�s%h���DI��;!�8~[m�z�[*k���ѩ����,a�F/�:����0���ܚ&(��H��9�r�]�!y��6;�l�ޫX�/1rz]����M�3xZ�>\I�D�W��������=�������7ذobp��M�x��ȓ���L_� �x}��}����vD���e��+v�;�|}č�z����K]ɍ��"'�#C��>|���fM��Sދ��ˎ�^e ��c֚�FYӑf�=�i�Bi�J�ϥ��g�g��>UE/� �73�2��րC�c��eR?��ʭ����:0� z�F�r�1cg��N���OWݘp�����V}»rw������Π�W�J�5O�.�$⿧A�
�D���J�(��P*c�|�����E�k�.�^���G@Cȧ!��n�p۰#t��[�h���ƹU���$-uL�����(��G�`���2���Ŧ^���w܂ĝ�-����3���j��{YwyU�#x���j	����l��Ͳ)-^����aֳ��YN�C_5w��GR?�D�j���1�M�_�v�� �`����L|��.�.sx�8p����Xeb����7��6/\����`������`����fVU�"��@��E�yq��啋�hʔ�]y���O@�|r�$2.#��}��N���5_�lZJH��7:��Cl��W��c1Z���H�0A��;�6�7���J�Ŗ���^�8K+���k���qx~�����f���q����jm�^k�����|�>��C`9s�����k�:!��ȏ��s�lgM��on?��x!3þ����<5JTF�U�m���6u��>�x#��i�֏E��2�M�BJ��l����6��SS� ���[m7I��0E�ۅ�Q0m�cs�gK���� ���F�3G�4㺍�M�l����%���^�掊�2?���/7_��&��9m���Y�D��g(�Ռ��w�c�l�f�f'2_�r�/gyp�ˮ��|�W�M�ΐS����w�U-�g�HW�۰����UӺ�ʩc��Z�s1�H@̉+W|�a�\	u���Ս�"�H�\AZ��Wd�
��0I3?�2��;Ke�
v0����c1��Kz��\�ޏZУ�!���B7d�sLEm!����hY���:���.��;����Js�%�'O1�Q[�'��˫�D )�#w�C����?,@X�B
�w�U�#�h�*Sa�)������#�zI�'������-��MP�p�>X���|���N�}�&��b�N�A9f��a��T�����cw�W�Q�V��M5����	Ko�A��Bbb�#i�;"ɺv��ժ��".�+�OA&��d�k��*�/�������C���b�lXdg8��īFjq-4,6��w�]����yf��]��m�5l�����V���$<��%�ΰ�G�[����B�^�]o�S�v�$Ai��2%��A2�r�#�KOF5�F�va�7�/�� �*[�N�M��(��iZ�>w�8|�W�4�����D �-�t���������GP/`lh����P���b��h�]_��̆|6��^}��*�2�W��	s�b��=��bqc��@�������b��s��<<��F1��q�`
`y�$>��c��[a ���f.l�g��y�wZ#��+���:��@7@�����L'u.��(ۃ����'7�)��W�@8����,n+/9��w!uPH`*v��̤�A������3	���+�[ՙه.Qs�tY��� ^[._��N������]t�V�k٠ث��<�o���WJ7v5;����ఞ��\{ؠ�3JAe�6	$x�%`����.���`�1�r(ڍ����(��!�+i�bmC��`�@�0�����Cm������%��L�g�H��t���e��E��~<�í(�y�r.A�Θ	r�Z�Z+X(��\�v
i�l{�SG-���-5����.!�F8ޮnJ��Zk�����z`鸫��Q�O4Z.`6e���5���v�n��k����=)�NtP��	.P�R�y\޾�R�&(ڦ̀�qn��Z��ȥ�Ja��K��W��v��I@f�w5��|rӍ�l���u��wV{X~�N���6ϛ3U���1����@9��NG���ٜЕZ������>���}s��r�H����X'?���w}'2*jo��'ՙ!�ݵ-��j���^fE$a�Ƈ4t�I��'i���/������M��?�>��_@��\�M��XĒؐil�L�ZQ6�ò���M-�XI�lL��r�F��#��A.0�:a��C���./lB�y��;�0��j��m�<��T��l*���{�~������mx���Se
�R^Ȑ�(D�fĕѝ�G`���>* �Z��VC�b�Y��E ��ՠ���P�FPD��{m����?�9�
��}27��gV�K�����v�����c<p[d0�V�T���t�Iv:C������%l!u[�N�۩����ʽ�@���"h�Y�t��K{�*zs�$�G�_��cÕ��F7[0zQHW�Q�e�)0�<9��	�Q�Pޡ����������q�5����NH���W���`IV��p�4Z�,:�a�Ch��%���o���e����"�^rc��󉀲YV���`g��/�)�.�,���"�s�H�����	S�|9�˕.|�Y�kOfb���r��ߥ�|�r�+e�����V���N�
�Py�H=y	V��p}�<-����o>�A���h�~ѫ������v�b��Ds�j�{
���"EZ�z�D���%���]X8T;���N�D�ى�?ӹ�u#��j��;�`BM�o��d5�?K��_���ΐ��Q����Sõ�񱚳��r*��#��+7��CL��g-���-�v�ݣ�(4Gzho��^32�r�j�hV�`}����猎p�+��L�w���1*(n�����5'���c���|_t;��`��+Y�I��9��6ڰ����`n��6lV,(.��y��=���[$1�!x�o�]�h�gΆ�ǰ�E�s��+�x�n�H���b|�I��)Ѱ�%�_ �������*{��V&Tl�$X���4���߆(��0;`�N_�"T�zL6��z���GQ�8?~fH�?o^�1��������D��guk8 V�*�
/z�7��HgS�-�P!	V��s&�GC�L����LER�����*�r��xlk8��rȕl��R�P��Ǉ<�5���m�H��7�)u#ע��[�B�9��K��/Ds�o0u!�R��I�K���A/�H��W��'����|?�˫��_�/��E�9��Ӄ���r͸�GZf|e�s.Lf%^���4
    ����          �  ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j����wEj�kB�A~r �x�2��H�"�BДN��á7ڴ �rA7Nm@��):Y�]��/�|��gW�:��Փ]���]�Wd���'��=�a0�a5k��7(��8�t9_����j�sRu�BMM�Dp��{?;b�)�����r/��F������Ό,�]��}��7�I�Ik�H\��Pnd���Y4l?���Y�E���Y�^�c(�w���T�w��>q1��/;� �#'o�Ĭ*�T:�(�^�e��\%Fɯ����[��� ?��`��<�������I̫-��(d:@��C'&é�1D�#)zL�Ԃ�/&F�}
��>o�x��I������k�aF�v����N5���Q7P��WS���}d��`��Y���ào����B���.[��8R1�	���q�q��m_D�Iu��8Kwݰ��Gt,D����$ ����\��R�E�o\�8�sGc�{8�%�2���{�����Tsr�lc2���G�d�I�a��G���Q5:�nj5_ٌ"pR]�-���J��xKÅ��@��"+cE)��T1�#G'r��b�SҘ3aumؓ��	I�Q��Ί��@��ή�%7����\>TE�?�S/���7ۍD����e�_ңe���j�!� ,'�t}�I��x�� /�� �6�48ݩ���&R8f�6�`�g!�4�_7�Rw�@a^�� {�7f.����z����)����4�&�G���Jz{�>����tU����Z��9Jj��Q/�m'�� #א���I&��>F���ڐ"V��[��Lڲ�02����؀���1X�Qw�4�ۊ�* ��A�^�4�.&�R��G�e��U�4ج��8DXD�#����3;V;��e;�����)G#pK%n��t7�ᔘ���O�XÇ�Ҹ��7�m��u`YӚD�y1Ü%��$6~�vKF|�9�x�9��4�Bj��1�j7O'*��1��j=��- _�Ԥ�p�{���g�]Q^q�S��I����s`��d���>���֏�a+���]�{�2e(��:l�RWE�����p&N�[H�
�V8�I$nť��b|������ 6�D����,A�3*�UXR��²O�_�ۇ�a\i"p��g�B����갦�����M3����)X1(����o)i��Hګ�Z�
4|���#Aj�n�?��<�jo��R���9yڽ�(��nS�ڧ%�ꪈk��8�R�-h�X{��,��^��%H峷�T��?���h"���3>����rx}�"඲�RE9�77(Kf�dr͛^�D�B�wkϱʊ!��T�kh��A��厚�(�Ӯ�.�P�������%��]����K�H�a���J��g#�X�4�JV�A���eg�n�.���lغ7��:w�''.��ΞU��o�p�N��XOQ?us���Ҭ<I�]���t�Cd���_Ca!k߿g�[���
��P;XL��b'f�m�ӄ������ު�]���c$�"��z4���x��{�V�
|�e=�ډ티��ة��F�f����|��	ze9��_Z�-���͂	�cC��>�F]T6�.���j��+��#Z���5Z�߇�MC-B���Ũ�SCL������ q����Oei��3S� R�t�d�%E�v���\�:ݒxl`���9��R:�U/ئ�0w}
�𠊠g:����3iTPn���r�RC�g�5=����n�>�^��lo�P��vA�� ������ƪ�6����E۩!�]{�u�����	�xHod�}*(����|�,���Ya84{�1v�sO���k����K�/���=���#&�;�6pKD�]�m0���m� ^��So��7;2O�����:�: �D��g����?_�e

���ysHUM�h�s��t�P��#y�ȁ~�d:�:�6LW��W=!��g!$�ϥ�/�o�����ɪ2�Xm�\�ʀ���Pm�\��zL�_}�/�+SRi[��� �
��k�gnt�)q��IK��X�
�2޵4��xj�.�p�
�l07 ��n	j�O^4ķ��������]�f��L�|��U&O��J���'�s7+��aO6N�=���#o��+�=!�y�"�p�.Y�z�;ф�h��J/.�q��ֳ{�<��}�o���6��>��fs	�wŴ)�&?�dk굜��xuL����ɹ��݅E�)鴿��a���HJ%RMW�ڴvV]m3	=�.\�$9�R��y�:��,��Z��7:K�m�Lc㮍��PQ*4i��M!"V�x8�FI�)ijWyv�'*.0?��G�f���f��0�21� �k(���!(��+�wp��u���p+��А�ρ0H8@�cR�&JY��ى�RO�Q�*���Y2.�� �VWm,i�o�J~Bcg�=۔n��+YR!"�aĤp�`��ޮF1�x�~Ϊ��N��R��0>U��b��g)tB�pe�d�҄cȜq�"��4��gC)��oiuC��&n�V���5pK��)W��Y�������~�1��fCђ�Zg#��[��u�+d{�[�,�R�=�X]2��g �=��%
&M/x�}7!�y�x. dߤKp���K�� ���c�YV�~��-дt�篷 ���r�>�C�-�i�6�Jȕe�`W!�������V'���{$��@����YB���
w�� �n����1{L"0f�b ��c6*���k%��s��l���o��?4�V��7}�|y���Q!(� �vC=��:U*��hzL�B���^ʓ���GǗ�\���{�pMC�;ec�h���
��Y��dh�������ږi���=�r��GW�Њ3�'pPpS�������2e������Gq["p��w>�N0��.1�C���)E����S� ���[�
L�$�]/�Qo���9�&Ke&Y@����4����8�,nv;�/<�=��eXt��m�Th�-cPs��˽�TKS�
�r�S4�-��6��ρ/n�`�X�cu�t�'�aN����.<D��)���� 3Y�>��RN�(�m��l��7P��#c��f��e���
�E�{}�o��U���*�?}�Y�����I����J�f:W ���(�U�σ�s��r@/�[�D�Ө��������Sأ�!	��5#�BkhֹhM
t��I#��h	@:�dn���_�� �](�pI=���K[D�ƹ�͌�IZ~�i�����4냼mm��PY̓���ѦL� ?UȦݓ��ۭ�(���q��h��
;ǥG�N �:���tY/3I�b�8����|/W�}K��]��vp?�$��U��Cb�Ϣ�]�c��	+�3��g�"�~c�p�R�k>�]�f��R=l��d�0O��/�����ECֽh[ۙ���H+�,��}"Nw)kKA�N�̝n�匦�S�U���@�Cz�eK�Zt�P�W8M��J�����I�?��I3����#�ܶg�r���l�N<O���K���}�΋�dF*�4|�5]�2q�%��gy�-8��Qİ���v�?�CA�$דH����N��kmc�@Ta��C�(��s `f��w��!��Ԟ N�r��3斲��#*Rκ
J��P�UۉR����<G��On��J>�xH�}��Wg|L.���v	���?�\�Eʒq�'�	��э,e���%���Գ�_s[�Q;�E�̴��o��Y�m?Ah\7p�Ո��O�B����Y��lW�,��l	k%����ї��JDF��-��[#����Q�2I�,WE~6E�/��H!G~� t����'aat�k��J�e�	rm�+��g3��c4S)�oZ8���Ũ$�o�Q��k󦝖����DST:�*m�_��di��_k�s���NL�1Ө�Æ׶��dl��w�O��i��jQ�K����Ia���$6D�;�O,d˼d�����da��n�ec~��D�����l)7��;��k��r�ԗ&᳃�P`��3�l�^o��6\K ��~��zܰ�$�V�=5c���\\R;�[�g�D�B��g�m�f.nc��z�5"=({&�����W��v&��L:���4�J ��?�O[+�%��l���ox����M����\ ռ��gd��JCt�Β����N�6'�]�w�'.�I!���աF��G'�m��O�Z����S�.�������ԃ:;��Kfp��"���C%�I��n��Ѿ�{� Ώ�7X3{��.4����G��4�6��#?�V���~��{�Rx�������a�R�īCq`�<Yҹ�k��1��t=���Y�"Y��F����WN�
Jf|�xW�������kke�<*&��b��;��3%���ڻ�:g`���9k���h��!Ӑ��ȫ�+G���"f �7!n2fQ)�݀�),��Z�-Ɲ���k�	 %-��X�'z��$S�iP?�w�·Ғ��z	���^�@�o�an�;��]S�������QP�YN���-��Y��n�z�G�%f��X�h�x�>�d�����Ւ����D�7�7^��PqҶ��
�Ot2�tQ��϶���i�	3o�P
�9״$�*{"�þy�Nh�tl>@��׼l
��bEln�e6"�g�/%�x>����<do�y`W�	C;%03�G��K#V�O��s�ۘ�4䪅3��|6x(��q��_��EZ�$&��6�染�{�MD��D���/�#�Jǆ�����.�F���e^	m&�,aPN\*������Gɴ�R���=44o)_o�
Gl�p"�<h�QvS?���*�L���̃��/DH	�L�\�i�_��=����rXX5U�ZՂ��X�B� [d��p��d<%���v����
����{�+�8#<�06h	p8�}��K{*���hsS��雉ܝ��s��������������Q�?���5�� 4:�u�=��Y��j���\����|�	��RԙW�M�4E���@�"c��>өd�*�C��l�4��d���^�d唫�E{�s�R���PI`�H͐��=��'��Ȁ02=m�,� �����Y�/f`g�ÃG3pL�^.�3�"�W5g�KItL����~Aq��{��M�бFg��{!���N�I�E$&��ȵ�~���y�����5&U[H�3x�"��V�d�o���u�c�l�dp��E��	�O�� ǂ� N�&3y5aȥ~ ҥ����' eC��J���ld"d�V�J��;<ܬc;�)���/����y�ܻ�s�ɰP��X�^�t�A�>P��%ǧЬr��l,;2R��ND�e�ܤL��ۣ�+y��Z����nR8&Nv��HS5�+ҹ�x�%�T��@D�_��,���Fv��Y�@	l)Y����nM� �g����Rm�0�R=�<(���$�D͊�Y+jS���e�Y����G)��je����n��\t��W ���Y%UD�� OFM�jk��Xf��и��'�FS���w�#�����ں�!s
��]3��'A`k89\ƭa��C�H������`�V�_X��3�[��ڿ���C���d����L�x���˼��ކ�̇�&)��[��6�o_�q����qcϦ��g��pO��-2ѤW��k���f�ּlCCN ��2�f�ݔC�����Α�R`2U�	��/��z�1�v�o���L뻡8��R���>%���i v�h8���H[��y�-���h���s���1���M�7�YH��2ӇH�O�zͺ�"���o��x��l����j�1��9�L�]���C�7��9_��Y��_q@:+j�G�*8ľ܄�����Q@^Huٌ�����Mg _��C8�q�X>LP�6z���1e��N�x�G|��8|���_VWF�K_��o�ś�惬�L\%d?�۰I~����!��1����T]u���I������D
H��z�^���&���,6��=�m�.0: u�k��o-�#���Y���	�?!~UP�)�ǜ�S�siM��-]R9��-��mV����Y�d�@(�"gR �7ǡ4h[l�L�����=Hk���h]�c����_��w�Z�+�5X_6h�X�o��!�2�Xg�^^͵!��F��ɔ�(�p1β�ܘ��,��7�CwNw$��0�ԓ���5�Y����g�l�	AU���4͊^��zL�����p�g�jlTa�t��5lP�H��*S�+�䁨��F��Ƌ��;�j u.��:�q xz��7��S��"�{H�V��l�?y_Ȃ)%�	�%�e���R��|,��~���������"QQ[JVP9z��Owp�g���+�I\�뇰�1	�Q��z��&L�,�Y���\�Yd򷦧6���kN�$���&k� ���nʨ[�zN�E�/�t��'7���(Y����-:�w$��s /
���5��7<�￪��o���I2Mj�����浥�_�)d_�g��)D�T���q���#_����S���(����m�1+4��(����?@�7$�	#G�M���$���U�5���k\�*�2�­���#��8JX|�G����;07���XF�0�H�Lt��0>	�k?[x�S�Z��bO\����aU]s.�],�2���lk�����[B�W�|s)��~��㪶Rw���{C=kB��FI)��L��)�M�T��1���Ztl��k*���-E&���Nkyyq����^�;�����.�P�����^U:���bG6O��������P�{iI4m���6Zi�k!1�uf���$�"��Z�;���h����F��u�DH���Sۄ?����,�@M�"*:�\��v���&�m�O���U�o_��Ϳ���(F��`�/F8�`NW��j����0c
��M�*����&����k�P����/�җ���ZT�7��AK/=��mnF�X����~��{4��=�}s��ݧ�g��i{�	��<�J?6U�е�E�99��tc<�� �B�<���k��/���R����Khl,�i��r�_\_%�4��R/s^Ȱ�`�Ρĝ�p9Q���^5@>oMS]��7G��E���zz�s�t@4�;}���Z��]�]�,[�k^�qW����<6F���*�mˤ B�ş���L�?�����E��9���~��~���N�j�c���]xVA��\* @����ۣ�g<M5Y��`���_��b�e&*=�}�V~��Q��B�Xki��!{sD�O�+�KuW�-�����r,��.��u���:�$d4n����\>�F7k�(�J�P������ ��?����B諔��ϩ�#��f�6yv��\��|��qֆ!?�|��_�E�/ȅ�Og�7�WGi5���뵦�+	{��zMϧ�^O����wې��;�>����l��Y�@E�`�/��"�zǍ� ���V��uI���˞�4��P�{�����A|ք����IC�*�~��2��f�ܥ;�6����$�K��#-x�a����y$D4a4b� ��s�+���ݲ4'��v�7{�>� ¹�hn�ƴ�Ь��TK�A�߶t6m,��&��@��V{:��Fs��Vv��%���
��̍<�J%cK#�;���a:o���Ի�Ź��`7��&��L��)�����1m7����:�Y�|��*EA�`Ǣ���*��eEX�$n��&X�����<�	Y�=�G��)s�6�)2�r�E�PDb�c��$���X䕵���t$��!o�);ǌH�
^��S���G�}xf+�ˊDd�q�N���F"���nK�4��<fCk��~I
�$$�xd�L1�
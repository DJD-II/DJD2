    ����            ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j�O�_�S��@�< IǕq��=��9WK1c��EK��ԣ����H�D.��	��T�����"O��#�WJe�l�Gxe}������!�Ea��X{�t>X��E�;E[F&����#�AY�����	�=�F�S�K7��i�ַP�;����Z�u��߮���S������P�ގ�D�D3R�3�����d�ր�^iD�zo�Xki��|�X"\g�}2�-����e����ѿ!�H����E{��d�a���H��AQ�����͘$��aC�-_moq��]\n+�����-�) �w�COdn�)���gHh�4�~�{7f�x0��.��G���SX6���Y�^d%<��t[5��sgn��	�o���>cj��9}Ր����f�R�����/^�f�.����Z�K�N����>-�?AäJ�[��9c��_@~&Gp(9��լ9ν|O���5tsަQ���^�$q!�)V:�{.�g�d��Db� �.�͂��4��� ����&r���Pi���V��;�|�
��������6�K�� t�P�TG����e��T��u�m�WO�|��_1k4�LI����,ZT�7E�C�k�s`Њ��u8�w�<n�,#��r���W���I���A���!i�!������T�Y$Rw�ĺ�T��c�mJ��oǽ~��ff�X�Q=vR���=K����k�T�>"|މ4�ܮ�5#�٘�F �00�ݝ�����1���*�m�*.*�*4�O��#[G�w���<��~�zUdM`�	CX����BlZ�i�ez}��=a��:RC�,��������Hh�k�n�<D�[3N�D��#W�EV ��e[mupL�j�;b��yH<����v��a9�������e*`���8��y	o�vΐM]�񳥪�`���^91����b}�8wZ�J�1
�k�q��z<�dtm������Qq�5wT��Q��)�Lң*�h%�4��
�_�e0e��(�U�k��P~":U�g��ag)o�L����m�`���Xt��mr�$��FJ�zUFȽ�ｙ��,�d���\��
N�i��e�����0U�ăX��a������.U��	$�A�[�*��c��RrF�^�p6�Z;��r��~�c�L}�)�8�s���d��ɦ�,`�&�ԪS.\xL���B�Բs��mﭔ�Mz�ʉ4�<�1`⠢k4B�ٹ�#D���n��lWB�|C;x�y��V&Y�
D�r	6l���g0Ss�s�$��<ĉ�z�rb_|���!�`��T�G5i�8Ī<
(+�E�,y%}:����p�Y��u����X
�Ӥ��1vP@P����������Q����q,��T�B-ޮI�)��<h�ǒ��w˒�s��h v�V&ssy����/��,�m��C�M���y��ɞd�Vg6ַj� \�� ��^�����5��N�l��(�q	J�N���i�|�J	�]vc �A�u�.WaX���z!���b1�A��H�-�xҕ6J�ܨ��N��3��qfP��#�_�@��~����)^��+r T�㤧"q��s4��#������Gۄ\��'��� ;����/���d�"�(��1ڸ���f�0�t����F���l������$h�E'�U[�.�J��Θ<���	���x����<rc rE:��CZj^!h�;\p
�9�X�j�~�s\�kR�����������x�e,�{Y*�n󃇯oH,��<B��M��< >JY5�*��3�g�����a��c}x��0��W�V�C�n�C3��|�8Am�*OQ����v���~檏9^Ǭ+0 ,�2��:��G�o��XJ_.�Y,� ��c����\%������^���dL2
�$�+m����69�@�<0�mP�[��!����_U��s�	b���t8�\u���󥐰k���B�<�kZb9����!�eQ
Cg��7�	Zi���0��m�6�޽p���4�s�`����#�p-h�D��/D
Tk����h#>���\�cT]pr�q.VW�H�!�!u�{ћ�{�ߗ�T�n@�#"���E�=Lh@�Pv��v��אY8���"���H:m���0$�����J�Z�UeKr�!�/k:&t�#�C�i�ˎ��7�,2�n[u׀�՛����؞�H������3g,f�#?Z����<6[߸&�a�{ot�A.�����I��B8�G[��'��u�����Uý<���;p��p.<����#�U]���o��5�S;�t�8d nI&N99��MhY<�Tc�]�y�T��N��Bn��<bڙ���\	ir&��94��7���x��7-�"YR܄xW�%P�y�8i�/QR��� w[�R	j&��ƙy�AD?�0�EFN�	�1����l���&a�Z� c3?���8�L�}L��B�xKU�������V���t���uݸK��=�w��4(RΉ$�^���撌����<�S�Y�Z^������%bOG���V�2�-�0-
��Z�������k7,�����ݐF�J�v-�}[� SO�@��V�#�dKt�^(��"��\��������8[#��v�x2ȫ���1�-8�$��;��Q��P6oO���F40�E�qI�^f�])�T���D��N)J�����ְ�4�]W��Ӱ���2���B͟^>�i/�ױ�l�	���QM[=$0q<��6%ՙ�ǂ���<��"�u�d#zV���t�S�|��r1�/���l(ޤ��$bkB��h5����˃��8,\��˱��r9���뛐��,)['��W3�)������� �b�Gf=����4|�&A�:�%I��|�G��p��2�'VT�qS����؅j�|M��RA�Y�{��>��%�u� wM=}����^ɧ���2�,�o��d3���k��6�/+�'�G?�ݝȅR�m�,ծ��Γ�0M�N���LF#��[c�5�e=Kmp�̑��FF���%Z/�Nc�zL/�1i �����3���s�T}2�������W"�e!2�6_�'[lbPSF����'�:t��Z�l�����w#A~;����N��fz����ӱ�>�vR�S�8�7l�TAז_�,�a2�e�v<@��)q��/^��l	mp#x	�µ��|k忰7n�ba3��(���_�H��Pqk�]�"Z�<�qu/.d�_�;�K�,\F(��^����t!ހ��8��b�+��σ��K�u�6#j`մS%@�t^�+	OFfˑ+V=�H����C�t���ri"�	��:p�����#D��վ����>����:i�������a����swGY�6���GM�Q'|�9��H�u�s�9X��uf�k|�8�b�Z��@���c����pw��f2r.��:H�+���LQ�drWU��2�*�9�"�I,0 (f�MB��ڪe��%�F���ݭ;�~JJ!�K갽���aM�'�;H�� ��+��7c��lD.,��r����v�L��Tv�Hq���������5�β�ek�S�VI~��?�q;D���Ս>��A�w{��C�R��2D�R�8"ͧ�q� 3�اPs!�����Iz���c}��3���)��a�#��"ڀ!��l�L%�a����^fAz\0UU��E�Xf"�^�j���/ftF�c�Vn�3*�蕭e6T��-P(yj�m�ZC٭�bo��UA%�YU$���3傃�J�����3&7t�˥�Q�B�� \�xA�W~��I�.�b�17HR���l���^i�Џ*���M3�\�/�����(������Qk>Yqx��w�R{'ҫt[Ŏ��N�$�0�� ���vP�"����Yw.�~n#��߽��-(�z����}fn�{��̰�V����Ս�p׈�H=�Ɩe��`�ئ�'�����(g�d,ꦺ�ԑRj�Z�����]%~�{.l��6]X��,w��f�G6�?T�g�䭂��Q.V��=*�8���8��I���ytj����
F����5����.����bM�n86W�2G�����uZ f�k>�6�"���TaL��2t� �T�+��:��@��T�\�;��?S�3j����U��k�M����&��uf�Y�/�����1�&(:�7����p�ν:�l�S4�1DB���u�b����_&�l{� � ��p�YL�\�6a�uhm�켒[td��LʲW&d~_��8�I���K����$ l���q�%CU(~M�!5K�_#�xR�/����&��0)T7��Wz;�g�7�0�J>�����>v�<�Y�G�؝��4zF�U��`B)+��Ͳm޴2n�bB�����q�f�<IS8���;)��/�:R��>�,�]�&�p7l,o(��G�F�E�y&����ᥖq�a8
T�KF�[��,n'hg����F��nRU��/�\k��y=p{�u�#J@��T_ޓE}�t��f��*H��f���*����zS8�ѝӗ�%�37���������z3���o������%c֦�Q&�H�pr������f"}��4��O��BUb��O�WkjB�|��o��$v�J����	�f���1pz�AUѾ�[V��F�F(se�vdܠvM�|o�%�����j�ű�V�̥g�|�/<���W�V��:�^���%E<��Em�.Y��������])`]��5p�I�]�^�'I�M�Vc]��������v
��'�R�����v��DHW4)5kà�S f[dI�P�y}������ǝ�$�!�j<o<�K�]�nw��(z^R��͵0��kG��s�U��i�Y�"����&xU�0���,\�诨�`��ǩ�;�N+*��֩s���k����O��&�M�Tc��\󩴛������ �$���W�!iοK �\�}z:�Ej�]�sD7j]psϔG9~��0u��JG��`5���7 a������	����x��xU�o�S����O*6����g�z���_�1L�Zq�|� 	�:�d����Ķ�w���ígR��.&�����>S6�ү<�yx1�qmv�����U���1?���Ma�X��tw�����Th�q�wB(�	!>��L%[zw��u��������䓔Q�tO��3�{)t^mb=�����l�����
͛�o��͗I��>p,�%�'�2���Xv�w��=6$GH�P-V�@)� QY�bݙ��'������߱A���������t�[E�Zw�]�Pc3}�|ߝ�M�?�D��&&�Kv�1j�N)�(�z7t�}
v���7�N}W!�@�2��j�r�ٶ6E��$"��9�w�A��!?Sm?"�!o�0d�/��X��@Ew|ს�u����[�"�[�Y��rf��.����?LA��'�]��;:>�"FR�x�\Rv"����'����{ïZ?��kߴ:���l�3l�wЪ}X��l ��-�a4������I����24�ON�p�I؂����m����*�۠K~b�\�F<��pʴs��LfO�X�8!�M����"�Aq����4�������o�	8���ϤE&ٶ����e�O{L��5�۴��i�mX��Q��ܦ�H��32�O5�]:��1Ϧ�����-�^���o��z,[�x�Ö��
?��i�l�7q�K�'��t�&��"Rr�+{���<
�	v�J"�3�γYv"��n}�VI�vKv9��X�
WdPo�F˨�5 �M�x�tr9R�����Qm�uF.���}n(Z�	M\(y28�*ȼ���d�U��vz�K�<�uΧe�"�I ؟<c�^ptm�q�j���}x�����w�i����f��o�8�{N�*arf+
�l��
���.�5e9�xRK!Nw!Td�2�o2���mq��q�	�_�r`D���-�>it�)qIq�|^�J��4���19,x�l�bIT5&�����P�'q�4>@5`�QBis7��S��p����o�O/�jP�L�c2����hI�s����F��D4��E
���d`/䀲Fj�쿹/����3�/�2�/���_V%�ldh�h�=A������_��:���{��0��P�
������{r(�����%�i�T{��',y��t�e�0��󕦹���U��TM���<��S��gIo��M�]��%�v�*�y���.���R (m�d@բ�3K��/N�*��+CǮVr�b�a<�h��/�I�Ʋ30:��A���&7D2��|�]��!|�F��A�"�~�p�תc2D7��%7�s�����9Ӭ��yB�`�W4�O��6�J
�x������T�A�:dG�u�����q���<��zp��o����05�5�{��Z'�)+���e��dZ_L�y�MR4�D�P�T�r��{5ҥ��ŗk��:�z��&R��$e��giƟ-��x�LX\�����2�<w	�K0�l�wM�L٘M ��r� ����5�������{%%�vZ�sʷ��rA-lE���m2[q L�7l�������Rd�u�@�٤ �$:	�������fry�L��/��d�Vs�쇮����tǁ	?{p�_�z)�����.�>�i��kd�ȕi���6'ew�,����3��T|�����CXj�B@`u�O�����^��� o���1��!�,�4�W$��Ż��T%��rx@�C�ftd4���a�����,{�gm�q���SI�ᘉ�=�?Vv�X!�`�K�_�/�x
=뀒I��@$�Cu�_9X�z����Ovn��Mǭ��0���hH)�[B�1I��!f}�n@I�����c��=����l�z���h�-罹7��8�Q4õ64���w{ء�?_$��@��*޷$��u�v��;��������;Y��s�־�v��~���R|J��ė��%м�� ��!�Ц��la��/_��TX�@�U!���E#P~��Tv�<��&�4?=�j(z�z"&��M1ш���+.�M��Rd;����~�6������!+/h&Tߑ��%�d��3��nI��<��j�d|��@s*Q)�L��'�öS�e���f2��M��7��� T��"~^�O�d�=,��%zq��	�;|�(婓���Z�;.���WX{-#/�H4U*��8�d�!-O@��B�j�
|���U;B��ddmN����Ɠ=�gan���4i�U�A,p�(	0!�;�)]��/�Fvѥ	�I���:"��]��Db?�ZA��~h08^��(��
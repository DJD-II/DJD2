    ����          �  ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j����wEj�kB�A~r �x�2��H�"�BДN��á7ڴ �rA7Nm@��):Y�]��/�|��gW�:��Փ]���]�Wd���'��=�a0�a5k��7(��8�t9_����j�sRu�BMM�Dp��{?;b�)�����r/��F������Ό,�]��}��7�I�Ik�H\��Pnd���Y4l?���Y�E���Y�^�c(�w���T�w��>q1��/;� �#'o�Ĭ*�T:�(�^�e��\%Fɯ����[��� ?��`��<�������I̫-��(d:@��C'&é�1D�#)zL�Ԃ�/&F�}
��>o�x��.����}����mW@�=����	h��EE���դ��H��"ّ�<5It·�9�U�s��T���$�#=�3ۤ��/�ʆ�����`�UO,�ğ������K[�i��C7��A
{�Ƥ��?� K������Ƃ�z�� ���"Q�&��QTa���d�.$6r�+��$c(�)$�����g�H����ޏd� ���y:E���}�O+�Q��X��;NhԹ���tƎh*�88�D���H�.���K���<z
lvmG,e�����7=��5鈮g�C�c;�O�,���=���2� �`��J�9���ȝǫ���Z�Hl�����v�ģՂ�O����lbg��E5E�����e"���P&���g��W��݇��,Jٔ�78�8m����� G�Wt��[^��� W�b#u#z��׈3�g�掵+ӻuQ������_�~��sV�'��� �\e$8#��c����f'iG
��l�����u�e6U��Лw�����9X���l���y�!����+���]��/휠t����:F{I|rX�� G#WP�X|^f/���������ir~vRZS2�����>�_&}�<{���JV��V��{~�:ƫ��t�!�qd�fck��<yh�l����XB|(�q����糛 ��[@��M��� [�':0i(ť�X�o�Q����Q��2P3�\����s�i-@5�9
,]�IrP,����W�����>�T�h�v�CK�L�o?U�����A�P���A�O&����s4�l��W�!� ��b-�ث�����B�T@��yB�ze8)ne��zF҉�M!�E!�<"�{��J4�FCm1�k��`U& ×4!^~�ળb�&�-b���*ʢ$N�k:���u��[�K��6C}}�����y˦�ֺ[�F)��$��1Gn�åα��T(^pT��b52�3������S�����@����'X/�<�:x�k2�D�z�k�'��\̥R��(��ZS]���ں��p�Vxc�U=�~U8<0�k�pF����Ո��/�q�lo��=[%2��V^���0��:d�	Ȇ+%�/�j������,2�w�@�!v��ϫ���5����������p�������J�*��N�H�CZ��TUR/�%�`Rp/���I�J�|\���*�4Ϧ�=\(���>{3`ѼpuAZ��3��T��E:2�4l�wwP�����I@�1S����b��V�y�2��G|~�w�9I��:����eY�巺S^�w�>[��>q��啝o$J��3�4��I��C�if'r
�u�I5��<�7�hL�I
�i�6�1j�~���R8��86MΎ/��M���z�\f�2�zN���S�1@��1$/R�5l���J����W4I�������1����eL5/���l�%Ԁ�Y��èS��U��hG���%Do�
�ߑ��h�Iʆ�C�61Fg�31M=��t��M��7C*�sN%��1�t�{J]�̓�˅��M� ժ����mi}3b+1ϵ��[-l2�@�YU�@|p��M� [Pi�����xP$�����WO<�%jg���HV��F�C��Lc5ׁkc['��ߠՍqu�Ա��38��0�*�ܒ�y%h���I<5�c�O����ހ����+>\�k\��P�1hs>'��0h�)	���[[5K�0�m��ٍ�!�4�Jf�d�;u�d6~�����0N�@X�3��\'���"G�6KL��s����Ѿ4&n�K�o��h*lY�e (�� ŭR��hD�f�a�l�����h��?l���A͵�{áF좰j��Gk� `0���!�V�H8q�_qL��E����)��¾��&=�O������?��vTa$ʧuFr��������������&^ �؞=$�+#���[W���$e��煥D��t�
�<��܈�����4��B=l�&�ڋ��z��'oY�����\���tmι˥T�8�M�at5���jc�YH�~.���A=wS�=P��^dGk��s3X-09��O~jT����y¹7�t�F�>�]���~��뫨y}��<�X�����S꤬��ZV.���o���h�P<�|���_B��L�܂�GS]�K��ה-���:��W�=���eȝ$�/�Ceu���u�`�6N�
��%?�/C���g�]i|*�ΈS)��y��I��������%��˝��wS��ZA���0�lA8�0׏kKr0�Ѣ�5���l5O��IX^���t'�V��o=t[�Ew8�؏�@�LصO���Z}^��L���Bxqȍ����q��s�������!%�}��X0 �6��!��C�IQ����N�k���71��Q؅�@Hm:@U�I�s)��a~ͧ�m�.;��TG�����`�ɫ�/��^�#�YhF@C�s�E��W 7}����<|�	���Ɵ Ϥn��&6��g��I�rS+���j+F��h�����,W��M���ό��*�`��b�ꆧw�,q+� i���+��|[��f��P���Uj5���B���13lnaE@�Xϔ\��U��k�b������0��!�<���,Ui����6�%FR�3|�ʽ�:�+|���ѷ[?+:���j^bv��<�)朰�����P*�=��5J�E!<ڈ���I�c �*T���ܭ4&�oe�S��'��#�$�Ӛ4Ep֨����Q[<[�4���!^����|n~h]��n���y�W�X���W��	s$�6X (U��>����)՟�rZ�jRc��B�k�0�N�O��5�m��sK=׾A��d7(j�9������	qAUT��z��x�I\p�aqf�/�F���Xxy�-Ѧ��ç����\]���ͨ�ހ��j����F�V��Hl�Z�p����\�Wr�D*���^���!n�oFLb�=k���\���I��i�^5t-h|vo%I�S�.ޔ�W��Ŵ�[ ��1�Z�NJW��S�s���W|����a�iY����M�q'��%�I�8��蘪A�`IEog3�Rg ���9��_>Xҋ8�Ph<]6
���>�s(K���\�:{�g�~��1W�QǪ�x���#���V�p�n�kB��-.��<r9ѬP��jL������q�5��,�uP�i�Qz\{���/K�@o[T�����ȣ�L3�"'J�C��8_����V�X�p��Ź^H�L~`{����:{XZ�'��$��7֖qz��Y��r}�с˺R��%!<��@�QR<�1�免���A�҆�_��z�L����T�S�.�Ak�m�g$#��޸�f	"��~/u=>����-�v�/v�r��!��;����,�6�����\60X	W�29,z��z"Oۨ$ƌ�ݩ�R#b�+���`�h��R;��-/|����O�8n���;%�5$�1���~F���!�H�\f͌��5Qdli��}�&��'�/�4�1.���Sqg�K�.)l���������~�([�h^�����<��vI�џ�1~�Py�r4A�%��F��o���19���#��X�Z0�Y�Jb�R���'P%�`!J�}���������W�X˲������)XQ�M+;�W7�tRØd'���ye���\�)!�-B�R<�>���A����ɕ0�f���T2Iik��H���E���C���'��̃�F�ث��2�y\A4��$f�f�t��Za.�&jr%��)�LS�����<g	-�I��W�n��%�6_�w�;|����'p�e�Ol��^T9�DE�_w:c��g̷.�}�f����\�l���T�79*1�/JE��qW���N範�Y��"x�%��j�	��0`�"f�tÛ�b�������d��c����HhbڒG��k�zBY��k_g�����e���ɪ1tE�o5ɕ�3)�ᝏF��#5��� 6�"B�l�N|5~�¤zS"�C`�
��1ސH!l�|&�apkl��i�ip����[�Gd�L;��6�7��Xh5Θ��b�v�����$p���MsJf�Y!�6��sdd�.p�����IW�[�-�03!����>�ҟ��<���}L�TÏ�#�S��;��S��cm�hi�'�����z��rA�����}��E��k6�)L�DdE0���I:D��ͪ�����c_*J����:C&��2c<��YN�4O�.�:n����\I# 4Y����q�N`m�ܞT�c/.����̜M�*��Q�[5�C����raq�����$���D�N2	�U����(���r� Mm2�}�������O��5yM�},�p'K��p��Pid�J��	��yF]Ut; hꦉ�7��&r'��5�-�d�j*��%ݍ� �fJ.�- i��a4�&���O��C�f��Gi�q�����>�m�syI�u+���YoPs�&:y�a�����9��^S�s,*`	�G�IZ	����F���~��r��}s��/fB*k�.�kV��]p�6SW���fކt5x<W3�5S&Z�������&y��g4��7d��bQ�db;G����^������;HhOut�jw��'ǐ�dP�ho�e��QТ�ĩ��RE��|��(a_Ԋ�i��M�� ��q�[����Ǜ���#[���pn
28KE�ʍM���ݳ�F$�1�PQ�>��>�HZ�h�0v*���g~�C!l�
Ȝ�VPM�S@����nD���ε`e�v�,�׼��wF�S~E&����$1��Z��B��u< ���J���6w��'¯��º�jZD	����B�v\����Ka�ʕ���}��q��ohE0g���B�
,�:ݢ����|ךi#�y7Ǡ����:�<� a�ot��3�,��uw�X�r��3s���CL�q"�m*��7��XO9͛;M����mb�����m��\-�
�.օ��P�A�n�����J8����/n��̜�)��)�/��}�E�l1����ٰ\�zs%l��H1��s���JX���q�|���B��C\�J�S�A����gK���P��01 �K�%W�����ٱd�S���S��i��7�^n�e�C�� K����.!*���_U��%�>��*�B�6��Ou�O�*����u���'��j�&�L�^�u��Ă��V��I��$���ѓ���ه��c����1QV�P��/0�у�I9�)��T��"a�{��������>�Zǈ@� X�":��@����&��Oi<�.�#Ο	/���Zg�Ť�C|�D���Z !ضI�ԫ����8��j{�/a�|���E��LlM$+�M���s+ͻ�8��{�F�JB���6F��_�dNщ4/�R� ��6ڳԌeh��@�̊$s`(����f���\u<�'�jG��t�Ɓ���?�/f���/H���":�P�qG����'�K�fJ�#j֍MNg��*�Bb�UVF�Y����!>��,�Շ*[n?�Ú�*&���_'s|�n���}E ���� P	$R�w��]��o��S���A�f2�c�F5U9�;���CC{�7�W�B��|b6�)2��|��U9Go�ܣ���{���'rB�b0%$�v�u������(R�.�H���y]1�яYdL*<��O?�b".� 
���nU�#��	Jە޷#mi�`?6v�4���RG�S���V�p�����2YU��S�N�k����)��o���ihnӻ��T=�"i���7�1��|�SX��3��l�`��N�@�3}4
���9&�.s�|�ӯiVI�����rn/@e=*֖ޅ\lN�tV!:Qҟח�66K��w��zd1�����%����GU��?B'��YY��	�����p��6�����ׅ�����E�v��L�Q���r4��OP�������󵸷rz�o��N���/�De��!dY[�G�x(=�v�Ѓ�fH�D���)]BE{�0~��=�	<��5x���IVǌkk�;�����$7��xv�N�q� eII��Z���|D���t����ê�ۗ�ս�S�!1�����J�=���聢����]j��a_vEf
��YءL� ���^`|�U������>�v�?���~BU��b�P�bp�J{�;��e�o���ઝ�l�ŗ}`;_���Mt�YO�G���T��p*EByB>Kv8�^��#�F��[kм�΅}�Tbn�5s�o��BK��(ӯnEڐ�o���+�r:ػ58�$���e�f%b����H�˽j��&{80p�/k�,�����)�v6���~��ª,�6%��1�f �9Քz����*�auB1qcY,F��������t��䶗��\��E&u�sV�#���=S;i�ǌ����¼��\h�Z����*Mdj�L`��ytDW�.�C
�L��Pvs�ii������?��8,�lW�&�n��=-�8��ȁVğ'���p�q��k����*������ͤ+S��ŻhᓥAP
C��D�(���$<8����r�Z����7�=n�J�������l{��3�4z<�w�/-M\.�8�ܙn�`�<�e�N�����]+}��&T�N�)q�a���{�w��י�L���uĈ�����53�2��~`כ.H>b��!{?��Yw���*�o�$U�櫞2��<.8��L˧�_�ͱ�cm!��]v^�A��Ww�u殨�^����|ju'��,9k��Q��W�mm��.{)����	���dh��<��m��ݰ���HF��d;W�Ds��QM�G%�sr{�8�AX�7>� ��;�f�]�~��O��F�=�M���_>(&k/v1���6����Lm��Bb(XЪ��m�p��(a\5L㬷���ER��9� �1`ib�2��͛���w6�B�Ig�%_8�s��7d>�.��k�b���D �Ƌ�K�
���艇0Q��j-�?ਅ�r1�v�L)֨�r�'�Ui��#Z�	����6+����W
Xm�Y)xP��v�JQ1խu�
_��x��!�~��Jɼ�]ח�ԋ;0���5����HQ%��4Xu|:�9^]��!I��}��0��;���q J���+�E2�f)� �"��C����9��W��O?ߪxϘ9�J&�����������gw�b��d��n���i;vt�y�蓄EZ-3��a�LXX�/�ȡ
�/�Z6KH�]�/�4P����������]f5M��o��_ȍ��'����j�"��`��'+# ℘.W�7�#�6�>mk��s]@�Ǒ�A־��Q{v����7��5�#)Z�xF���(�_T��Z��}��B�_��"v�[��p)�]W��U��&I�( �Jt�6�Y��@g��j�7�#$i�Zc�.��p k��v��<i]Щ�7Gj�DE�	N�rrF�taI��7���o�Mue��G��>^y�����SO3����q0�_�x�a\a� ���0
s���Q�������/�(�o��֭k{�Nw=��F�JB,Lp��O��j��J�t��#X�)GE��%�7f&�
    ����          �  ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j����wEj�kB�A~r �x�2��H�"�BДN��á7ڴ �rA7Nm@��):Y�]��/�|��gW�:��Փ]���]�Wd���'��=�a0�a5k��7(��8�t9_����j�sRu�BMM�Dp��{?;b�)�����r/��F������Ό,�]��}��7�I�Ik�H\��Pnd���Y4l?���Y�E���Y�^�c(�w���T�w��>q1��/;� �#'o�Ĭ*�T:�(�^�e��\%Fɯ����[��� ?��`��<�������I̫-��(d:@��C'&é�1D�#)zL�Ԃ�/&F�}
��>o�x�ۊK�0�M��P�hH]e�� N}��#e|�ey���.����g�Xt���Q�E�r�築a9�$������u�w����:u�G��Z\P l�/��9-ng<,y�Q'�|�b��(�ZO�@��W�Get0�T_�|��ѰZ
�� ��&��	�q,(F�p���M\ޠ��q�!�3���P2֏��{Ĕ��K��G���>�O`��U��*��{Wo��� K�ipDB��I7
͝����>�K��� ؞}(R��c�(�����jw�4����i�im���!s小L��j~��7!����YG��\�R��f掓$~�E��h���~��Z���{~(�Ί�n��5�~���D��@���"��0��Lg%�fjiAs�%��n���ay�{�}X�q\��xb�cʾ&��)B[U'�1)=�T�I	$\a�����"˙u~��T{�$��i��V���O�K|mHt�[e��)P���2�I��Ǔ�6���)�����=�#VQ�� �[}��)���NDmhU�ZJ�{倿Bo�L��6�"O4�*��΋x���IJ>,W��YП��̇��+I�0H�q�cۦh���y�:x��{�K��8u�FT�+D�M�,��<�{4;Z�����3_�WT��/vl�X7.�J���$l]=�1��o{@5
X���{P�ky��"έ,�W�w��K�NI+2����:�����9�6�иe�W�&ú%�{�6��L�_!�=Q�r���S}�Ǵ�� <Q�妢�r����K���.i��������l`�޵zg�@��	�j��u^gQ�_�O�"L�o���)����,�j,�8?�tp��)�O�Ҽ��Mi�_,]i!}Y%�Nu~�24�����4��w\�W[����f���xOL0,���`�y��*g�?۴GA�B�	s��Y-����*_n��?�ҞNPx��B�φ���%x�Lqv��N�Vn^3n�,���l���k�"H�l�KuUl{7c>�|����S�]H3���8t�����R�J������H/$���҇�CkJ��������Ùܽx�1��5ٮ�X�c�
�xVZl�r�l	J���d┬�j�!9���_���k3�j�6�a�Lv����E�G�����ʍ?,(dnu��Z!�T��gm˼拔���&�� e'V�V;�>�A.����|��I�V�L�� �FD�`�ab�l�0���5r.q/��?X�n��Fɂ��梩B����d�w��)��׋UA�
;׻S��B6����9���^�P�:Z]2���!�h�^T�я8��Ls�ټI}�<?���["_"���6G.�'����Foe{��YK��踏��4��>\�lt&��b�]��:�RZ��;Q�Jr-� ��G/_m�m�|4d��Н[_���	>��Ũèn�����Q �,�N�p\���a�#�m�+����&���sZ�j_�e���W��-Z+*��	���e�����j��f=�+�^#�H�zY��24})��M��Ұv�t�)�pY�� ���LS�48w~x{\:�fǨ�:0�	��hvDK���m
P�qزC%w�!_�QI��HO���	�H���m|�g�{+9���Q�ޢ�$�R�^��d����?�X#��8�ǉ\�VD��"����k�nCB`\�H�����y��$�@�N����S�!c�����Ml�s/�e%S�l2���TT�񉁩��(��"�^=u�5S�1ڃ��� Yw�+C�C����cTC";���)1aol�z���P�z����f>'@\������ep�@�?wƫ�3�@P$���|!>��m��dOH5'e��4$F��q6x�q��4��R[�Y�R���M���8%�<A�<5IOk�B��_Xn��!�����X��l ��|�"#*�Z�()�WY2�.��$�����A�w����^4(W_M�9���TR<N�'����y���mM�YH"dQYg�8u���[."�&TAW�$��`Ċ�ry��� �r<��U����_\�RIО������VLl�lt=zT�j�KΫa� �+��C,���*�O{<�(�Ō`�Au�����܀w��:�܏�;��BԂ$���A�yF���t+j��H0��9[r��^�O4�4����CC$�6)ߛ����y�M]��]�>�t�߯�	�	x��͛7m>�gu�;zo��2!��Y���3�c��9TK
V�ᘦ�*���G�|*H��6㖗�I1�мv�<_iz[%���ڕBz$O����˗+^b9�9��:L�=�H����1��-I��@'�ރ�^i�$��b�!(*��	���L�60K���2xy����������+�a���j�����Oc�d���#�з9�r2���F�����O�U��Hs�7y�w���u
����Vb���p���U�(�#Ǘh�PU��߽�[B	���l�� +��yx���9�
�Q!QM~��zG����Cl$������t ���%���)��z	��
�@�k��������ʇ3쀤����.��ݵ7�.,�t�Y�s-^Fܠ͝k2uI��^O�I��zo��[�As@���1L@�v����k
t���W�u�jFP���=)�g�a��I/_��\�M5Ҕ��������"x���Z6lP�rL��s%��1��n��)V�
����m��q|�����雩���`9#��]i����	Z3a2�P!�2�_p���y�ӫ��LX�2eo�!�����l��Ii:[��r�����`��]�Y�	����]e|]b�t�!�
���3�&Z2��<��2O�x��I㵐��J�`Q�������E<m��k2{�Ȅ������,�M��{k��z�l�D=�o%`�g���F	���S�P2`�"���a���Ì�?��ܿ���ȅ����W�`��3�3��^����,D�,?�"������`��c�z�
����9��
�i�sVƱ�7�Ȅ�ö�j0K˕y%��&���wO��NKh�ɲm�WضSP�q�k8�E�y�<*V�`�O*ocq�ft�����y���8g�-� U����{�I�n�VK��m*�P�ϥ�}�y�Mdߗ����(8(����pW�e�=R�g<x#��~F��,9�]r*�`K㕘�f��.��i #�!�h�'��ɤ�3�o6ڽ���#�WB9��h�kR�߁)7��yeiv~����#Uq@ܐ�5�?��t�������H�\��V�פyp�?Zf��'#��mx��!��Nu՛��ϔ{5*S��ob�vfZ�k�B%/>u/+ʗ߅����䲡5_�p�˰B���E�@оt������,�ekX��@�9������"�܏9u��vN�͐�߃�o��]�0R$����67¡J���fۋ�@��;�q�}�G~'|�J)Ϣ��	jR�+��O����8�f����d�EW��Q��ݙi�)r�AB�#?��I]^W2��%N��h����a?5\�I��kn�,�%���:� G�TՈ1�{�d�AR��	�$f�Q�2i��f��_������Ѕ�Z�m�6�ug%�l*?(H+x�H�>2yD�`�RQ�ci2�A*�>�Q�6v��<����=����B�Ϲ1�G�搵��ٟ���=P��P	AK@�T��>H>7�Ac�1s��k�9Y�	2��h�7r#� ����}��1�ɝ�D�u���H׉d�o�{oL)/��JCl�L���=���+ aR�а��4�v�]%'[ʺ��F��X:����' �%�8��5�Ft#[��l'�k��
=Z(���i	�rP:�vR��[/���a�χЭ*TuV,�/֥�a�i���B�����X8�4���?���8!O��
���Y�y�j�ǟ;��W\���i���f18�ʵ#Sm��;�Δ�j��)Eh=�
=�H�\R�̉U-b�WO^�v�*2��%�Hl��$��Gz�}�o9^�SJVܴ���u����������7�`)6��~;ij��7����uŃSc�uWfw�>3ZxFC�}-��[T���9B��4�D�;�{M�5�]AA�-��è���?���9�ʇ����Vc����g����gY�~�)骇8ϱ�jE_o�X3
r9���m�>ːY�8�U�(�ln=�+��Ӻ[�+ �l�2��e��PQ�6����!���H�[�IR��j��xm1�&�Ϯ-yP�D��]���7(dR�C?w0im���e!(�h�* �6|9ۈ� �F����.�����
'��|�9%�gB�d��J��DdvV����'���F��Gز~�4�}�`#5d�U�mMc6v���QG����S$}�!�)7�le�=O��$H�� ˁλ��k}���]�(�N�ak�/2)��A}�]j�P]��HƂt�������.��;�Xz=�}I{7��#*��g1�=|�+D���v_;�F��rR���!S�!�?mtC���Uj|�$��j���y6|V���5j���x�C���'��0��7���|��h�Ҕ��М�vmFL�&�x��Yj�n �Ӂ�C���TS����#�K#���I���o>����S�N����q�җvj7; Tf;�^�����F�9籊�����?�S�ݾ��?c� ��}��А��c|�l���|��S�S�(.ø�}q���񸞳C�;'�DV�n�n�\ׄ��BY�[Mk+��t���QS�T���\( u/�i4n�`]�ChL��ԏ�i�t?z����y�����^�~j�w˜�(���A����YݕK
	;�RY���A�#@ܯ`��~�n�Ic�B��X7�8���g�ƙ���8{ l�`E�X4Ř<ӗ�U)�����D�c��]ޒ��+�aYm_dhE>�O�Y��&��m;��LE��Yn��_W���2����Z��Wct���hΙ��ؾ�NN��?)��i��#ȦRT��M��y�eR}t��Ư!�9|�1Z7��ϴ��	=_5�6���_���׬�ߞ�E��|�)'�+�x��u$'탔j�ǋb�H7Я�ؙ��K��Di���ڍ���z7i�P�B�(�R{N|�$\��AW���r�����b�N�L)c6�^@�ߒ]���,����-;�͡�﯋��<{�{8ecn��9`Wo����M���A�H��6f-�:�s�ܕ�L���9�m�Vsb)i��(�5������ݼZ�� H/6Z�w��>nZ}t�@}8�q^v�4㬋��Q�i���:�<�Y��<��Q��Bj�g��f_/N�~�y'���q���	�29"�KwN6���(I��I�����­\M��?��C�C	h{�Ҙd����3.
������x�\�qp =�~���)l��6��󶨌���PВ��)}Q 0:�(��M��~'��ࡉ_a=�m���3$f�&��a(XӐ�	}��q����]�>����Sz��l���*	*D�J5�V���K3�s�W�O��u�R�w��'j��n9@X������=���O��V5e�����*�B�
e�b�6r�Oj�'��j���h�V�eN��>��9Cc~z��v����Q 2�.O�=�N���q����麎{�y#�>s�V�|��P�{�?{Z���v��=�`X�#�u{�f+&�x��6ng��F����������&�G	�$ЊR��'��e�C?��F;��S�	�hA,y:nm�a>��4��2*GϦ\Z K�]m&����m_m������u��D*�٬%�*},�踟�P6��*�T���*G���l�f2��@�Қ8v��?�������(h+0R#�|��45�j�'3 J�5,I�N�֞���WT;=2�K:G}̆d���mb7�\�����_J�\L�#������_�Q2[s	ರ�s�#\I>˳�Q�b��`�Zߵ��I2�T��M�	����K�0[�r��)ۏ����������6D[^7�[Z�t..�M(�����X(���Oo�
	��ᙡk�6(U����xY��,Cvb|��9-���]�����g��De�)��Z��D0��W���Q:�a���Z���̹#=��$��h��_�u���E9����8�7�,@����۠�KV� �6�X1��tb��-��ŧ�&'��<�B�j�"������噽k�#�0t�$BĠyK~��c��s";��a(��TE_>)61Zetqz�B��;�@R�jSǈ�<�����M�;>.<�`����#|V��(b�O����E�F���I�y>7`�Yp��1��8^ͭV���GL�lx?�z��I�"AM5������A��3�	���`\��'G�(�UlM]3��-����}Q	6f3�W�#F�M>s��b���lX��G�C�����2]_�����Q,�6�Cu �܉�wb�[��;�|�O�	�{�\O?��Z�������48�1ӫH��H^����I�/���@�~SD����=�*�Ȗ32X�Nu��?<�{t�ǰ��ۄ�i���=��ML 굵�-Nю~<�܍�w��0��ڛ��RO�I4 �Z6G�1�u���Ո4�Qs��R]\��:������7��9���.���X��*��lZ�q`�.�rÏ?Kg%.�-�^\j�}�7�:�2�Y�� ��������p�����*Ҍ�t��1�m+Tcl��z]X�VE�E�ဟ�d��e�����r�'���a�;ğ�OꊻPi�`EmE,����6N]���J����>�C�-��a2�55���O��l ͏Hs�`ײ�fw�XU�ȍ0�V��hޅWy�;�i���H�i7�m3����ٕ�줪�fȳ�=�m}�C=�8O��1��Mht\Þ�K���)�N�r�L��£�T��̏,R�qe�o8l���	��gK�����6o�C�2���> _2|�~��..����Ew|	��fHR�_�����Lw�!�dC9袟	��IS@��5����m��\���u���R��>B�� 6�l��u�&
О���µ��6F�W�'ґ���A�c�z$�l2$+ϐ�9�OK�ɼ��A~��{���W������6}/����*ZW��sn�t��E��D�^�xP��aL֤Q��ȋ�t8fnD��Wd-c�F\rƷ�-��4(Yf�l�i8�貱�φ�篝h�~��G�L�1���CP5�+r��
f�kQ���/,r�%�m]��iϙ�����!Q�����L��s�w��vO=j�L'��2aC�|�⍞��%��`���ȼ���������FHq�۞��8y~/�M2�2���]�@�y��,Y���Y�ͷ��$�uX�b%+�ך�7��x�	�a�F�p��+R���l�th͋I��c�L<�A��R=��c�)�Q�j^l҉�6��e#iG�7�mO��.�_*bc����v��F�^}@�A������}Ա������Ʉ��^��w�\>Oå�o:�ʪ
    ����          �  ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j����wEj�kB�A~r �x�2��H�"�BДN��á7ڴ �rA7Nm@��):Y�]��/�|��gW�:��Փ]���]�Wd���'��=�a0�a5k��7(��8�t9_����j�sRu�BMM�Dp��{?;b�)�����r/��F������Ό,�]��}��7�I�Ik�H\��Pnd���Y4l?���Y�E���Y�^�c(�w���T�w��>q1��/;� �#'o�Ĭ*�T:�(�^�e��\%Fɯ����[��� ?��`��<�������I̫-��(d:@��C'&é�1D�#)zL�Ԃ�/&F�}
��>o�x��&�ٖ��P| @�$ܕ_�ܘ��r(�n�ٖ�����Δ��O�6*�B��^�,}�Y�U�$eg Z�C�Ys=ܯ+��r��2��T0]2o��i��
�(d�e��J���W���C�lR&��.�Kv6����_�bY�|�� *��d��/���U[��+��p���tsg�3S��*s�c�R
}��}Y�G+ ���Z�S���+�bjN�Y�$W,�����	Ԭ�2��V��{�e3�h���~���#Q�3�Wj�|��H��`�1��u�j:~E�m/g8H����S���Q�|MΜm����_6Q�~ :3p���|�N��uB��R
��*y�UO>5=PISL�rE�P����BX"x�����U�?c��/�z�H
�[����M���Y�^3����\X/Y��������4�[�`,���A~EL�]���v���#�4Bs2�B��n,���Z<���5�̡�q��O��x-q��ZOI��,�{Mv����y 8��煴m��CwQ�73��ݬBx%���8�ڀ ρ�*�D���}�D����u���C�(��G
�pe�A\<η�#��oR����Ҁ��CPV�ѕ��(�!G�򨱦��O�y���҃�������X��?A/�Wz����Un�����ق�f����_˃��c�T���t`|���]���J�����<�6&K��;�Q2h
{|_�3�컫W������s� �y~�T�y��h7�ԝʪ�<�x�m�pG)��:�*��${�DY��T���<�}`U�K⮔�s�%�ߙ�a¦֬�٫K���,F�D%�0�bH5�ɀ}wg�Wf�n�́;P(��1,��j9���+[4)�ny�}f����͟�U�W\�K�-��;�kbp�9/W�z���U�E=�#�FS>O߉�~�;��40H|Õݪ�}��n|Ԣ̛�]Lf	v�OpY7�d��Gk0\�.O1ؠ���X����`�K��|��>����t�z�?{D�>s�R<�C/P?}�H�h�{G�b�M~�IŢr㝙�Jz�ZAn[ q�$�I����hC�B�(;G,��L�Nv\fr�29O�֡����w�<S~�^�0�l�	��@���$������Of�I�c�$����'�\��U�������X�!����sQQ�*
!M��6n�X�o�.�(G`ނ��a���\q�hH��W���匊��JfM�Q0RY5�֗"�����Գ���:��\���y���0��4G����"ؤ$�	<��\����W�P�N�J��Z�qL�1B1�	x�,�����W��A�+��q V�p�=+|��fnC�p#�G\�{�n�X���Iv��/�4����J����o�R�ۦ^��˳�LB6���zCu��ؖ��̰��V]|-o�;ߣ�m�`Yc�����K/�y��,{��Gi��Y�P�7���iEt>���!xܓ����U�-2r��P2R��~��x[kjO���ط'�Z���P�5�W6�=)�^��ʄO}i�l�Z���&�"�R�-�T�q)�Y���;Փ�4�٨G�:-��1��j��V���\o���GO ���ʆ:��@��0�:�����2�8Z��޽�"�.��G�Z�QZKp�-d��_nL�Ȳ�����W_��4�U�?0���?���4L+cOM&j�-��$F�L�Ý����VlOZ�}TF�6�X7Y���3�j(����H��9צ���Niw3�� ;nVxH�)Ҽ�\�������|/�]8��a���s�3�|݃� �	eZ�M=�-�����4�6��rg��i�,-6���P���K�y�Uͷ,�_�\���>�	����vN��ŷTo5��yBx��XO[�7/5�e��PO�ьE{>���v!��Jg�fQtZ��	�>���"R3��&��I޻}"���:B?�d��Ea����������]�3����ZD�]P������\'��\�|��j�yz�Q���(���Ͱ������ /�ā�fL�0�h3D؏������L��؃�-uv�Y�p�ޟϲ���r�qS<�5�����j�P������If!21��  ��BtA
P�x>b>Si�v�}s�i���s���\E�AO�5�O�Xb�ޔJ���go�R<
�"���?��B9���2��p��	$�6)k�V�ut�h��<�èHO�i��� ���^~��}A�~�:~ͷ�[ci����`���[Ȁ��to�{6N
h���p!�����ϛH�ټ�֤IS�{1�����E����&�T���l���%�G�#'��J�yU��|eӍ=晨p�uG-Baɲ#L��#�Yu�;�=��H	Φ�����,a"��7���B�ї[p&Om��(π����~����.0,8�Gt'nyNk��4o��V��ɮ4���O����r|882\��{`f;�6��]'M���k�ѧ�f`P[�h�\u�4�g�w����:�U�!y��<پ�ՙ�T����=��5����Muʞ��z�	uQ����ɳ�w���/ų��m�&�A>���(��\T����V�}������g�����eIEV@�KHzh(���Q��Ԇ
���3�z��XPx����~�gw��1t6�,�:s�_(��d�3!��&<�ͫ=�A�|3�knt�1ǥ�hg�t��R���ǛZrƈaZ~���X�lYcs�W�,b��f#V��Y�_��P)��4�&�X�{��rBD
8m�i���.d��"���@��0�s�
:}���~��@TH��_����A�.�B��n�u������Mѡ� #�����p�#�8�7��~�i�1�B~I辉0>\��.�U?�����'�P�R �3���ܤ���/\u�:�,�B�1uh���������w�Y����㰎���\�|���������?>1zw<�Ђ�:%kbof6�����=�Z�&	�%WO�X��"���F�K�) ��{Uܵ�ڞ��jqӐ<��ע��JC
4���#���7�-W���Oj����S�WIyiKL�y���]}�fc&�$�lR���[��C
??�$�@I�#A�a���D�����G6�Ck��%SNGc}+r�DJh��v"�Q������6����g�*5�y�M�dKҖuCj�\�;P� ���I����M�O(9�k��e�N? �g�'�=z��RU��{p�{h��@�7���J�V/���ؠD�k	�#6��>	�P^X�:�C�~�ò�k]�%~o*i���t4��(��r_#��&qr!�q�̿,,��鼅2v���l��~_���U�%��#l��aJ־(�\�8�=[�~=�W\)NBoN�L��	VoV�'�t1=�a�0�8��!/Gr#���H�[�NR�}B	�*|%Q���W�Ȼ��k�_y��^��-�
��e��p�s(6��Jf��(h�9��8�Kq�_�{d/�����y��1�����#uY�eκ)�8i Ns�� �ߋ+��v�rQy!��곦3��!ܥ>�>�;�~���Z��x�gh�A�}q������!PTY 7k�/�f`��R#\r��w�s�f�r�,ǳ�ny���$�w�O��J�y4��k��G�����j(ݞ�<���zg�A�㩳���7�3�nq�C��G����1�x,Wc*�.~���V�,óv�x���2R[��$�ί�{�@��+
� ���5��F��X��Gx��.��<�cM�zc�;��X�ND!��=L3l����y��V7����x,1Omt�BGq��F�{*�A~4Q���̄gC��T�a}�y|76=�#&�S>�����G)�S����&.Z��/ݺ�t�]Q��9�6y䔞c�ѣd&��z:SDB%I ��T��r�M�|�	N�*��2?�$���n"H� 4�ሼo�"(I�2��A����̡CQ �|�Ԅ�{ٲp�à�<�1�����%I��L��;�G�`� _��1����˸��̶�>�:o�\ ������O�փʹ"P|���N���U��M����͋��mW���#��9��pJnr&W�cOt�w'�RQyCg��;.O{KB�V��T�2сqR�HT�'��i݋7�W�pDեO3#��3���S>�]`p���8&k�L��zw���qi'\ �j�kɘ���װ��#I=�	��0L.�-K�d�G�ɡ���`ܹ��Q	Eˋ�v\6����0�s|��z�9�N#͍�/!����az8�M�. �+�s-0�¬��&�����ď�d@t�����:��Z��J@І�z
9��h+����ۄʷ ���i��w�r�g4	w��;����]}ky�Z�:h+�z�a����&F���!�E4sE4V�,�S>�0�3�X��4�,f��(cޙLJ��W���,��.
�O���1^�D�F�$M��f�7D�"�½�\<�0ʩ�ʀ�m�g�D
�d�:⻰钚��3�Cgpי!�䂂,��k�Q p]11�࿏���1���
ؓ��o	�8f?��k�������`�Ҭ�W�ٯ��wF�����i/d��J�2�6*�9t|���.OKK�*��d}P�����Q%�����_·�Û��#�\HX��A�5���8韣��oTw���4A�
zl�j�\����3X�/58��B.$��2H�gDP�A��)q����f�T:�t�'�&���+�s�� ���Dg]�Y|��̠��:�I�6ZZ��A�Q�s{����F�P���d�íd�/���.Bo�n��Ŀ��8�%a�\�IW���@i��"9��\ca|�5s\۔����	X~����g��x��`��k@��Mq�Jz�9��L���+�)���:0�5[���g����#� �nH�`��o#���[����$u��WJ�R͓�D�cX+�#�~m�e|�7��/���|��>+��i��\=1��Du���ԅ����v��2�;�`(�HQ��siԜ��=��>A��8��ʲ�Jz���Z�V۬�'ć�O�\�W��6��t�ք-S-���xn����;:�;����ύ����i浚\ͨ2U��h��{��4��=U�����Y+>�1e~O$-��Sz��V�t�E�:���uw�%�eg��BLMtmϔ��R:O"u�h��MJQVtO��K**��"�DmRG �u�7�g��ʢ
f*~-k����`�a�%b�q�5DU�w�V9>4TT���\�����>�ҹR�VB�$�Z����;��u�R��t�n�o��_�T����K}�#�=���:�R�����3���,��ޙ�d����0����W���CmY���m>�ݚ�"��:�槔oq�PWɸx4�%bW��������fG�-Ig˪(�a�#z�C�v�3�c���ÀH>��{�@CF�y��k��I[��m�{�i�T�V�,D9� H-֟��>@��6ߗ��Qs6S��6M��`��V�a%�̧}`�:x��Ku��@����<^���'���5g}�i�_�wi���Э�JI׬NUn�L�v�Д���K[���d��׽��uBK�SF�g��#Gm�]/�Ex�*�{7K����r�#���H�|��p��|��6t�[aR�ą��K*�>�lb�ʂ�5��u�>��[�G*�f{����2*��Z�|��MM֣� �eM1O�DM�[���$/�BlB��/��'{�2��u'7�ڊ�����N0�]��j�����h�%,�x'��Z�/���r�5�t�`�������lZ������Tz#��ޛ�ۏ������ߟ���>�C^{dy�^s˨�LgvCP_헠�a�O���5�mmk-C����L�o$�8�P�7 	��������"����FHF�X��k�f!Z�������f�^Zá�x~x���[~l�Q��Ŭq��j�B����R������I�Y�e��!��+��~���
4�m��Z�Ę��q
1QO/+��<@oo�{LX��G~���wLMk3O��_A�r�L�t[�I��­�z��4���������;Y���H���v��u��������l����X���"	�>��N��ު�'���OA3f���Ƶ��X�|�-�}H*"D��ME!��`�������;2,Kɸ�ft?����;Ch_����sC���=�c�ײ~G$c���dbUc|��SA%ZW��yj����k� &�ܘޔ	},$~:�)JA���O�tR��tm4�pz����)���}F3��Ї�pp��d�1�?��᣿��\����~�+-g�7�f�"�k?`�C�S�m"��)�Q��'?����K�Up�8�_y�Y:�^����������xTYfſ-s{�����_--@T�niZ,��9ul�ד��m/�ʽ�(����S�f,N�o$�e�}6�����.�5@f�>Q%UΥG!O�_1�o��^	6��>��� �C��W繅ӧ�ri�?<���h=�nKHL@l�.
�?�i���f6�݊O�VR�%�_|-���θ���u j�+��_�_����~r/ �*)�"�%c�hOԻ=��&��g�v�>^e]Ep.cJ�2K��l'�*�lW]LK+҉0��.~��yMZ �����	������է��uJ��g����_ ��-����!i���@�A��M�����t���'a �����s�R@��4�����ûF9��S�y��F/`�h$��)<r�^���tj�&y��b��( M������+�+\�:�ػ>���/IB�~v7��yJ�}�$h��N��Hk�ʉс$iW1W_���~�!�P��X���2Y��d�z�O������=��v�c(T���0�c^����P�?\o݌�W'HK?����ș�.q���|��Z�.��E;�>>�Ĕb��,�,�F-���ҏ��jv�چ�&z��0$n��T��A�3�I���m(�>t�k��K:��Ѯ#����w&�0��{�KL�ȝ��u��+��_ ��������1u���y��Ȳ����˩Y@S��P�
�<�TA�c��|��.u�Ĉ��Gv��2���\S�T=�W�a>�u,[��|�U˧����@SGT�)4qF�LlE+ۚC�^�c��F��*O�O��ǃ|P��\v�f�X�3���g����Q����� ���V����s��/��?&~s
�c0��@0C�s���h*B<��D^K�{�����"G���r}��|c�جUU�
��׏N��.�/S�!�S@�QZP����c�G�(
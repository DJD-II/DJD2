    ����          �  ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j����wEj�kB�A~r �x�2��H�"�BДN��á7ڴ �rA7Nm@��):Y�]��/�|��gW�:��Փ]���]�Wd���'��=�a0�a5k��7(��8�t9_����j�sRu�BMM�Dp��{?;b�)�����r/��F������Ό,�]��}��7�I�Ik�H\��Pnd���Y4l?���Y�E���Y�^�c(�w���T�w��>q1��/;� �#'o�Ĭ*�T:�(�^�e��\%Fɯ����[��� ?��`��<�������I̫-��(d:@��C'&é�1D�#)zL�Ԃ�/&F�}
��>o�x��&�ٖ��P| @�$ܕ_�ܘ��r(�n�ٖ�����Δ��O�6*�B��^�,}�Y�U�$eg Z�C�Ys=ܯ+��r��2��T0]2o��i��
�(d�e��J���W���C�lR&��.�Kv6����_�bY�|�� *��d��/���U[��+��p���tsg�3S��*s�c�R
}��}Y�G+ ���Z�S���+�bjN�Y�$W,�����	Ԭ�2��V��{�e3�h���~���#Q�3�Wj�|��H��`�1��u�j:~E�m/g8H����S���Q��(m��%t�H�� ?��������av5�>.:_^�ⳡ��0�^DaCZ�T��R&��B�Lj���j3MU�P���W7��P|��]4>��]��5�|1<G��ͧ"I�|�^|<����0\�}m?��dIg�4�wz a�[1���)Wn�'5�]��n!��h_�K{��U��{�1iLp�զЋ2w�R��0TB�Tm� �����3�ӭb��iBb�,�}�5J�V�'�S�l⃧����!��*ُ!��{���ÿ�[�.�n��˓з�H�k�s��R�H�Eߢ��M�sSP@�G �âi~/SZ�,����?P)0�KO�
���3'����{PΣ�˾�������V�?���L�jsͪ��x`[�c��N�6�� E"�n%a��<킔y�������[���z����J�J�8r�/��c�B�K�%�����N�m�A������P�u1񃱗JQ��Gv���U`�e(u."8��ۚG��7�c�@�92����Cu�7Ը�"��p�Wm����]J�,��W���)ܶD��#�
P�U�a}�{���A(�Ɠ���W�"�U-�z͊n�S�K~W�hM���J�0��]��e���{��"�(��i�M�J�0����㥱m�\=Q���lBT��=�&3�nn9��4�Ud�ms����:�����ǘL�U��ƚ}�Z�P�|~������M0�R���C�A���ߦ�=�f�E��c/X��0���>�s���`�@J��KD��{vi	�ʼp�ӒWȏقd��eIr��B,����6�"leXk(E��.IC�k֭�mi��`�i�Y�;g�LA��h�ۜf�v��늻L0�b��[#퉾��	(dyْ8����"�2л��%���y���W*� 8���QF.��)lr ������n�-���7!T8����7c:a>���oh����Ө@��B��s`6l+�غ)^���#ڏ<
����������f,/�f�D?c��K_|Q&�儔|���H����0���ř�BÎ�'��e�B6DA<9 �p7�X���l���+/��"�y�]:�=@�����w}x�m1i�BMZ���(6�l�
,t?�W���=O]Y�;��uدF���R���N�5��+�W3�r�},ZF����> s���~K]=rk�*���K����ʆ�^w|�����2���-���`�uz��9������x��O,I:$t��n�I鵟޻�0��_�u��)��l{����g��kn��<95�A�=#7#��+��m��@j��$G[8QTB�5ގ����
�B���1��I��j�߀�8�8��2�y��A¸��5�X��	����8 &���F��yT�i"�Vڳ���0�d�H�Gl��e�a�d�W��yͺ\Ղ�Ѹ߮�8r�{Z��cӨo���k�L�J8&�P5�&ݔ�o>ߝ�|�~ڌ�A�m��)a��׵Ke%�����5�]/\�ܐ��x񒖥׼«�hPuq̽�-��7�4F6�����Wg�ߚz���w�N9Y\���������*0�_D�z���ޓ��x�?ɒ�@�m�_2���\>�w����	�L3t���P�M��y[��[@%�uc y�s!�<[�۞��pXN�cHi��=c[6Y��P�þ:=� F��`��th6�Or`�}ʊY*��p;@1��Z�.�ş��z=7M�v;e�����3o�����^y���+oN��`/��O�`�Mƴ���L ��ƾ�{�M���A�$pؔ5�����u8G#C���(��m�s:|x��=[���_��"�c���B����mhW4��K�9�Pk��k�/*r�4�)�͞�r�~/ǰ&J���0�hk���Ak
��G�+��z�������zL�L#��%K�K׼����/Y.�D������`�km_k����e��M&,T?X�+l6� �"��{~�ǰ���8���č��qV�.v���Н��l�c��R�����\>ܼzV��Ȯ���Ɓӗ���#��%��^{n�r��n�2d��q��7"b�I�s��y�M�<Z?���ĔQ�b$s!��ͧ�r,7o۩k������9�ɃT�^��Y��`��7�| 1�����3�V���X�"�]�A�]ŘBV�)��*n׵�5�}����W�l1iЉ\���6<G����hui��P�(1]�A��O�c~xe��۾Gr~y�:-e=��9��[m�%b��Q�:i����+�uKl	�&��@��~`y�~��7K�Y�ĮY*�����p}7
�MV�$�������6uC���������5!擰[)�E�#�9(h�C9{�2�5�W�^�{rf+�w�M�5��B�o��!�e�ފ�B�暻�J�h���}ð����G=Cv�U�E"�|�xC8;�^%hXA���G/���W�3�6����0�(��U	�+or�צ�T`'_��:�	U���@#����+B�hk�c�9���	\�͠ɬmP/b�s.t���	�vlr<-��椺�)���L4��A%�Eo(݈�1�QI'Z��κ1�� 1vC�E��f�6 �F�
Ӿ�ax9��w��ꉃ��սr�,M~|Y�h�9�g���z�/��:��m�y�����Af�-B��l���e����������b�-ҧ';U��5���YAn:1N�H��|zE��#1����Sk<�@�w��`�]V��:z-�Cof��`�jטe�{�=������?��?x��ymk�x$t ���c�n���n�n����\}څ�� 4��������Z	�f��K�����m̋�{c�&���b:�|E��-C��Ͷ&f�).�]��]�/��R�e�^_����OԄx��J�ںA���C؟ό�D�ݑSf1R�s*�0�g�l_J��-���a�8C [H���9=|G�:�+Z-�z���O���r"��k�'���M��@G|���sx"H�bБ:6-n�����6}$%~o�!н�Y���X+[���7R%�W@������!��lȕ�NxtD�u
U�W�AF�q�vvb%���> "�i��<�B[�A>i�'���gTK����*�#u�Y>�lV����0�/饗	�9�㚞y��qb�e���*�uT�nw�ƛbc���C`�0���;��p"?\z�!ZN���m�v�D��Ym��	;��GD;��C��9�Jކ�
�B`"}z�t�~][]�i��n=�p�Ǧ(�`�I_�!�(*W�ʊw�UH��	���G�ox�66�lae�1��<4�Ƒ"{߃Oe�S�0� ��V�gU���@T ��^H�InBV�fԿN9��b1��5�L5w�E1�N�$�� /�<����{���7�v�G�̪��
k5|Nw�C3�)�s�Y8	q�{�i!��p�J1�����e��M�y��#�&'�q���H ���;��g=6%\g0���e���'�=c�I�71=}�:"��)�`�S��޾��Ye���
F\t�Vk�ݶ���@��'d�J�kT̛hx�k��+��̺� 	�8n��*-(?
��}�s�������A$�PE��cV��ի��gB4M��`ۢ]���6㦐�0�/]�4�[T:�⼪�<]�:��',V��^�B�K�.���� ��Wfo@@g��sh5"Jc,B/�K�Pt����:���5�o���=�'u@s9���%�|�ZR��	c�Ƅo���L�^�=^Z1�k`#�������^�>��ӯP����r ��OU+����+cH�}������땎�¥+� �w{�Sӝ�N*��%�'�3��;����|e+�{.��K�l��wxp��#&��ӘM@!�zm��(�$#�q!��s�"ۍw���wtc�$V�:VM�P|�3n��\4#�?uR-HY�dorÕEգ�]��)�pw�VV�B���֮���� ��pC_�w�R��]�]�ҭ��m �`���U0ro_�F�{8�I�C���>q��e�˸�Z-	J`Y� "?e"�exx�f�[�g�4,�bR`"'�Xa���A�����$'Goy����[����v��i�E�I!Kd)l��+���v�6��ٚhבK�����������������w�cm]���>cQ?iL��� ZQap/��o�z L]'����T���
�^��p���>����?�s��_\[���t-ɒme@�l��^H!aKB���Z.�8N���`��8N�lw<�LC�%o�#gm!�z-L ���O<����>?��L,�99�T(�DK~C:ŝ�M"�7<Hd�BmO�'�a�����ۉ��N>EidAi��|�W�U�\H
�1"'g@��C��Ք��/̝�ŝ����gC��{mn��k�(�<�S���a��Z4p&7��^���A�+���3�mU%?�|�}6�����ղ��|��{�[`�UvM�%��ӕ�ߞ=��rX��r�� ��yٞPƵp�{�Y�%6a�}G0�ZƧM�32���y��?�?�r��y[�ރq�Qd��r�>l^����[p��0�%H�M݅��C�Շ��m9!�EJ �K���ʛ�'�?t�^�17��	=���0f]�)O�k�\��D>����y!�w�^)rAw��)�N c���ˑ����%3_3��$����eL�v*`�ܼv;��֠f�����w����Jə{�
K��"q=f��Z�}-B�aݚ4?�~�ͻ����.P�<>�q�P�K�l8����i`�3 �䉓�i�CF�꾡">\�`S�}��څ�ῳ��H�p5w�o]7�d�tdp%�ԅ�儦ߜ?�SA�AX�j�����˦�M����.2�+W��6��!�|8�&=D�HpΝ1�[���߈]�+2sk�k�(x�0�<���AIJ3��?B�؅6�-�`�P�RD}�ݨ'!@�z�(2��J��e�
���J��u2�E���XG����Q,��`�ɉ_T �2���9���S-���[����Z�N��+;�@�.C��%�g�rB?���!՛k�c	A�G���Rj�d(��%O���p����cS;�uUa��Y@�r���Tm.)@9X��L�Y�t�_7�3���ڰ�D��%/�y�VH�s�"�,���_U���ȑ�� |h�P��L��]a�����*U�;lJ�@_D��%��!DId�AXoK?�q��G����}��GWA���a�Q����5 ���KE�<�tW�<�w_yI�\��e��̅�6���F�z
?N��	�jz"[o�L���O��?1~O�(S$�$�~�d���N3R���JڪXɅ�~pJ�z�"������l��2F�.<KEe���+��y9���8|�Ce�?��� �n���l����E�GN�h��=���-�6��3�&P��R�L��?2�)`9�Mj�Χ_���Y3�{}Ϥ�]}|���<����N|!W<���r��U/C�T_�����a- �/{�*c��hR�]O�5B ?��Q㵋ˠ( ��V�#��|�U�,�zw����x̨�z~�^%7o�g��C�`���E��Oځ8�F�qJ��S%�;L����7���D�՜��'&oD���]�-x�΃F�]Nب!%%q� ~E���L&�s�1�%��
�gI� �pr6jo�p�y#�ӄ�S}�`�N�4���G�V����ҌX�d��y �f�A'��/ϛ�P�C ��׺T�BO�wWn�cI��]�� \��W����F��[e�.����}��%4w�u±�Di����s��`J��	�k�͇�#/�Q:r�4 �0=�rTa8���(�vH����V�?jT���UMY/Ó<�F�5i�ʆ�b��Q�ҹ6�s��Q���8rpm�+()w���*�Y�gs9����!��)�|��eo�'l�ȯ�]=�>��jۑ!���d�����<^��#O�eJ��X�K�2K;w%��:��Py��L������
G5]m��f��iK���(�:!r�4ll������{�?�Lġ!!��Q�����/��B�]�C'�1�!Z�饔}@ٵ�+��\㊶���kJ���o�kD����7r�9@^U��^�n�d7ظX�f���t�������M\��*'�r��������V��#^^���T���e����d���d�#�?1����X��՚������ϩ��������)��B�1�3���Y{֟o�ʹ7�I�ܳ�<���5<��ҍD�<<���OE��$m�6+e�&�����:�����)����#�V��Z����G�I�G���"��"���R��a�}^��9!}S͂u/��������u�1��v�}G^��P�*Q��YQH�溧@� �!���3&�Kv�㆘ަU��T��0�50@��� �i	�� !�� �:b=v�$�V5n�x1�J5-w+�����/�)6F�?sN��d�
늴�O�b����0����7�SY����/�(�,��8?b
R)@N�$�J�B۸���S�+d������$~9ِ&H�w�+��4`�w�9�t�P*S1��>E��C�FGl���:�ˈ5jܠO}r]�fa�����[��zm�������p�>�l�_�y�Ã��"��O+P�r��['�]5��u��\~�ĔE����\���3ud~��?�?��Ԙ�����ı|MR�2bl����s?�1�H|U[����&���v�Od�m0�}��+³-�Sd\�'.�/xO^�G7T����
�T������rĄ�֏��w��H�
��J��9�<��׏s^P�}���l1I�יP��*�P�txs��Η��\����9�����J-�KG�IiĨ
�M�8��5�e*�£.�Y�
c֠'��&��Ƅ��:�<ng/U:���������c��e�mw{�:2�����[ï��B��v<��d��b+�z��t�	�(�{��@am�=������ߍ�Q�{��R���IrrЛb��ķ�"��{�U=� �͗����|P��q�o���"�3T빾s`�V�p�5����Sdi�.TĹ�P��\-c��L�R�X��vBæ��d&�7A�� })&w�]�e�7��n`�GD�;tQH�u���\����z0B9�^���z�͈Q�+M7��>t�ҭ�2�H���%�S抳}�Ě��$Mq6;?��_�~��O:WýϠ���`����H���yX[�<�޴
    ����          �  ۧ[�/��'ti�í|��O8�Ye�dr�#7z�ל����WUC��@0�PlD\�g߂η:�O3Y%�
�?Φ��\i(vB��XG��D�=f�t��j����wEj�kB�A~r �x�2��H�"�BДN��á7ڴ �rA7Nm@��):Y�]��/�|��gW�:��Փ]���]�Wd���'��=�a0�a5k��7(��8�t9_����j�sRu�BMM�Dp��{?;b�)�����r/��F������Ό,�]��}��7�I�Ik�H\��Pnd���Y4l?���Y�E���Y�^�c(�w���T�w��>q1��/;� �#'o�Ĭ*�T:�(�^�e��\%Fɯ����[��� ?��`��<�������I̫-��(d:@��C'&é�1D�#)zL�Ԃ�/&F�}
��>o�x��&�ٖ��P| @�$ܕ_�ܘ��r(�n�ٖ�����Δ��O�6*�B��^�,}�Y�U�$eg Z�C�Ys=ܯ+��r��2��T0]2o��i��
�(d�e��J���W���C�lR&��.�Kv6����_�bY�|�� *��d��/���U[��+��p���tsg�3S��*s�c�R
}��}Y�G+ ���Z�S���+�bjN�Y�$W,�����	Ԭ�2��V��{�e3�h���~���#Q�3�Wj�|��H��`�1��u�j:~E�m/g8H����S���Q��(m��%t�H�� ?��������av5�>.:_^�ⳡ��0�^DaCZ�T��R&��B�Lj���j3MU�P���W7��P|��]4>��]��5�|1<G��ͧ"I�|�^|<����0\�}m?��dIg�4�wz a�[1���)Wn�'5�]��n!��h_�K{��U��{�1iLp�զЋ2w�R��0TB�Tm� �����3�ӭb��iBb�,�}�5J�V�'�S�l⃧����!��*ُ!��{���ÿ�[�.�n��˓з�H�k�s��R�H�Eߢ��M�sSP@�G �âi~/SZ�,����?P)0�KO�
���3'����{PΣ�˾�������V�?���L�jsͪ��x`[�c��N�6�� E"�n%a��<킔y�������[���z����J�J�8r�/��c�B�K�%�����N�m�A������P�u1񃱗JQ��Gv���U`�e(u."8��ۚG��7�c�@�92����Cu�7Ը�"��p�Wm����]J�,��W���)ܶD��#�
P�U�a}�{���A(�Ɠ���W�"�U-�z͊n�S�K~W�hM���J�0��]��e���{��"�(��i�M�J�0����㥱m�\=Q���lBT��=�&3�nn9��4�Ud�ms����:�����ǘL�U��ƚ}�Z�P�|~������M0�R���C�A���ߦ�=�f�E��c/X��0���>�s���`�@J��KD��{vi	�ʼp�ӒWȏقd��eIr��B,����6�"leXk(E��.IC�k֭�mi��`�i�Y�;g�LA��h�ۜf�v��늻L0�b��[#퉾��	(dyْ8����"�2л��%���y���W*� 8���QF.��)lr ������n�-���7!T8����7c:a>���oh����Ө@��B��s`6l+�غ)^���#ڏ<
����������f,/�f�D?c��K_|Q&�儔|���H����0���ř�BÎ�'��e�B6DA<9 �p7�X���l���+/��"�y�]:�=@�����w}x�m1i�BMZ���(6�l�
,t?�W���=O]Y�;��uدF���R���N�5��+�W3�r�},ZF����> s���~K]=rk�*���K����ʆ�^w|�����2���-���`�uz��9������x��O,I:$t��n�I鵟޻�0��_�u��)��l{����g��kn��<95�A�=#7#��+��m��@j��$G[8QTB�5ގ����
�B���1��I��j�߀�8�8��2�y��A¸��5�X��	����8 &���F��yT�i"�Vڳ���0�d�H�Gl��e�a�d�W��yͺ\Ղ�Ѹ߮�8r�{Z��cӨo���k�L�J8&�P5�&ݔ�o>ߝ�|�~ڌ�A�m��)a��׵Ke%�����5�]/\�ܐ��x񒖥׼«�hPuq̽�-��7�4F6�����Wg�ߚz���w�N9Y\���������*0�_D�z���ޓ��x�?ɒ�@�m�_2���\>�w����	�L3t���P�M��y[��[@%�uc y�s!�<[�۞��pXN�cHi��=c[6Y��P�þ:=� F��`��th6�Or`�}ʊY*��p;@1��Z�.�ş��z=7M�v;e�����3o�����^y���+oN��`/��O�`�Mƴ���L ��ƾ�{�M���A�$pؔ5�����u8G#C���(��m�s:|x��=[���_��"�c���B����mhW4��K�9�Pk��k�/*r�4�)�͞�r�~/ǰ&J���0�hk���Ak
��G�+��z�������zL�L#��%K�K׼����/Y.�D������`�km_k����e��M&,T?X�+l6� �"��{~�ǰ���8���č��qV�.v���Н��l�c��R�����\>ܼzV��Ȯ���Ɓӗ���#��%��^{n�r��n�2d��q��7"b�I�s��y�M�<Z?���ĔQ�b$s!��ͧ�r,7o۩k������9�ɃT�^��Y��`��7�| 1�����3�V���X�"�]�A�]ŘBV�)��*n׵�5�}����W�l1iЉ\���6<G����hui��P�(1]�A��O�c~xe��۾Gr~y�:-e=��9��[m�%b��Q�:i����+�uKl	�&��@��~`y�~��7K�Y�ĮY*�����p}7
�MV�$�������6uC���������5!擰[)�E�#�9(h�C9{�2�5�W�^�{rf+�w�M�5��B�o��!�e�ފ�B�暻�J�h���}ð����G=Cv�U�E"�|�xC8;�^%hXA���G/���W�3�6����0�(��U	�+or�צ�T`'_��:�	U���@#����+B�hk�c�9���	\�͠ɬmP/b�s.t���	�vlr<-��椺�)���L4��A%�Eo(݈�1�QI'Z��κ1�� 1vC�E��f�6 �F�
Ӿ�ax9��w��ꉃ��սr�,M~|Y�h�9�g���z�/��:��m�y�����Af�-B��l���e����������b�-ҧ';U��5���YAn:1N�H��|zE��#1����Sk<�@�w��`�]V��:z-�Cof��`�jטe�{�=������?��?x��ymk�x$t ���c�n���n�n����\}څ�� 4��������Z	�f��K�����m̋�{c�&���b:�|E��-C��Ͷ&f�).�]��]�/��R�e�^_����OԄx��J�ںA���C؟ό�D�ݑSf1R�s*�0�g�l_J��-���a�8C [H���9=|G�:�+Z-�z���O���r"��k�'���M��@G|���sx"H�bБ:6-n�����6}$%~o�!н�Y���X+[���7R%�W@������!��lȕ�NxtD�u
U�W�AF�q�vvb%���> "�i��<�B[�A>i�'���gTK����*�#u�Y>�lV����0�/饗	�9�㚞y��qb�e���*�uT�nw�ƛbc���C`�0��^ݝE���e���=����
�R_�3 �ܤ)�y\&պ{j8����Tc3�~{y���hE2��@������xYvb��H�[�m��������2��{�G��G�7����Xɰ$�X>�S�0��E�ba�E� �M�}��j(4j�hK ���p�%�Ka����>f��
�3�aY�B1y&�#�|�o�O��Q'�Ο��[T8�l���}�x6�����Q y,z��V�� l����>+2�@ƚ4��#�**>�қ,�2�Q�X������ܧ9u�N���5ƩQ��V�T�=C��$���#�0w�{����K0u�\ؐ5N3_����Msa e�UCU��%��a8�i��ݖA�2�uMP�t��C����Y8�H�R)x��n��J�۔/�e���9`�d�	�Xa%BF�C�q"�'̊�с�����6���L8���,Mn.O;q�ٯ|�����v����,�sDтT�YX{Pm�X\�h!�M.I�^	��!�A�3�5�D���'�3����T�}�.��%	�Q?�l��
�Ylt��{6�� �菷���|�Fa��ԃmMW�Qd;�(��(W؆�!q��}x��FY�kQaB�t��m����+��]�h1���%ߪj��1��(2�������t�����C�~u����&�~�����(�Gf����(`Lh�<3�n�>�ϥUݤM�K�8�=}��mbEZ�jÏ�&�4��,04ʄ�'�6��\,�)���k����!
���1�}ڕ�D�Al��lBX��#Oj���}#L9�w��K �W�Q��[�	Oio�3��$�Qv�*��v]�<�o����a:}*�5o�E���C��mC�xkY�7kKM�w�c�b����XW���$�㎋
{3�44x�����yk�E��IN�K�(�$��9�Ҿ�<2q�2�cXTs
>��1V�?�>�K/���
z:q�69.h��A�w��P���hI��3�A��u9�Oh�X~|؄B&"�=���O~�i7Ù�������o�ZM����x5R�W��GJ#���^����>a�O0REƜv.��|$�$��xF�4`���03�uU����� ~�����lh"-C�3������ϧL������c������l�U}iQ{j�h	�i�.gIm� ���I����ɂ��1BaO�g�P�#_�{�4n���U���ƒy����Bf��v3$�hߋ�=a��L�gG�~Ғք���=�(Q{T;�.s׃����G��a�z��WJ�ʚ�zo�Ow��B�/�8� ����:�/�C����8�V���D6�n뽮r��D`�7�Ň��o�X}ߋ���Kr��-	�.l&٦�-::丒�C��od�Q �X�}�sp6�H,J)��=|l�������We~5�v� Ih�?�����3|�J�Q�v�VՃҙX񑂚.��p,�6����]Aڭ鲢>����W)sm[_�N;
)��xHxB2��Z���Q�UQ�m�>���|�_3�$E�'y?)¤�k��C�'��# �;�d�jO�.���ca��S?9!�+����Q�g�֗S�??L�[mڈhuz&�����ק��W�6A��)���J#1[3���s��-��\#��>$A�<��j��Kie���_�w�`�K�f2���٢~��j�926�fGTt�(�р	��<�Uq����@ 9���4W�1�O ���'T�N�Uc��A���x$�l]�.�.����ڸ�7W�"�A��Ӎ����h�A��a3��?ػ$�R����4�7�՘��Dڃ���j��|!Wit��7��#*X�օ�P�*h�_L_�Ơ:JL}V|��Y�Hs����>��1��u���:,���F�,�E)ձ�V�����j���Q�*C����d-�����#�q�n��<��?�����b<``p��x��2ؤ$	�-k���>}إ�5�ב�V��	�Yr���jMȸI�F!s�1��;�1��(}�Й�Wc8h�x�qM��D�F�'�o�(��nk��cm�E&,�El��C�<P����R���+��|�ے.X��mhNh���rUIh0��TMd~ڑ04�ؤ��&�{��u�Ħc�ѺޒEj�Avf���V�
�� ]z��Od �:d���>������!-Q�1�\&��6�+��2D�3���#{ݞ�avW?����o�5�3��R�Q�x�0���`�d&���I�7�zx��!=蓹��H�u�V�ŉ.� ���h�W�J�Q���5B]�~o�+sM��Jd�k��foř�j��'�.����dW�"��\���|j1��$����*�����
�f`{ '~���~���)vC|ͩ�4�7��� �C�1������+���jK �tDp�w�XX����4z�P�y��g�jQjƦ��uH?�f��	�$X[WQ}G���k��@x�y���0������O���[R�I��Sd�o6[!L�NX��[^�}�!;�6�{��n;p�NNf6�$\�	�d�&��Q�5����FW��G �e��M�&|��8��>�h	(�c�krĩ�f�?Y9�|g_�x=�X;v��ٲ�tJ}��������X��=�l콠�5ck����Ep	?��-	;��] .��c�|q�o���(�������'��y{�/�{0t�K�'~�z��m""0�Z��$��N8@vǹ���x�H!��S��I��>�XSp��Iа�h7�Y���)�]&�}��>�P*�Q�P�h�P4f�f+?7���o�3��)7����M���\��ҷ���Hi��1,�{��G����T'���.bAhBa.ݪk�3� �c��HL�s_��˶,�A�%vBI���)Oy��η�kG�x��"/�kF�w��r�Y��t��<c�{��ِ�<����	?�(����'�T���D����@���ȅH�ݞ^
Sˉ��˨��2�@{*�������f��M��Q&vEH_4�,��?-4p9̢� ��=t�d�x��Ǝ��Ő�o���`W��.�Gb�wu��`P���d�;! �8�8.3!�]��G'�y�NCb�`�O3�o5��zo�l<�u��|�h	1��c�B�)`/Җ!-fu���D��g	Jr�𹔣`!~�=wF~PR�2�����Ж��V��v�H�@�_��/�&�J`ck���:�9lU�W���b+���_����2����* u�� �у�옰`�&\
��]1� >������ �V�λk�U����ړB��YawK��NP��:<��h\-#�IA�|��oW�-DJ�:i�{��R��w�9[ʠ�ۦʟ����w�ZD�]���""d�kvP>���P ?��jʸtva�ޭ4��A%�!O7�mdR'�0��'2����[X���CǾ+0�t��RU��I���7r�������ͩ:P_ݗl<��n��	x0_-�Ҩ��~���:[Fx$9=�>�PƼ��7��#kaڑ4�030WU۝0w�Hʵ5���0����_.��y:#��K:J����F���f�W��>|�KU�1�]G~�+���I��cx�c�6�w�Ͽ����ۆT�!�����^9^�.���T��O��1�ʊBȗf"�@j��V��K=���ø\O'��� O��`m��ZW��2�<��	?�#M��IH��&O�Fڵ<9u�G=W�H��,��Q�C����ޓt��+�/S�Ro
@�>��O�d=;�*T�	���T�"��Z:�u+��42q9�:��>�l1���V��'X����H�K�_��앫\���I-���Q������,(�
�g%�'%b}B&�>�rb@K�k�͎/�E;n��SXݨ��s)��tr��El2+��)���h�|����W�	�Π�FI��Q��[������ۍJe��q�^$��U���ߪ�3��a��qs7�����a�C�>�:�@�(��	3�0fz��śA���x����je�kX3�I�'9�٠� Vl��@��ad
�h�5"�e�����S�`�A�
��������mh�5�f>	�RZ�#źՋ-Y��_bn_��a)}��"��|k��ơ_C���;_gAk�t"�E